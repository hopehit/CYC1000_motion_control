// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:30:26 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MTLMq79ip+jLp7sp6SyJgzSJ3KuQzDoHYxwFFpdt6re7oCLX++/rKVGrTpkuYpZK
XNIAFVmvk4QZ1wzCLkCSATEh/kpVlXeEX8iiew5Rrjl0kX+xekfpM6LXnN4fLnfB
M3T4eZgVoDfjM2AW058mdr9d9vLwYV70BXHeAErLE5s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33584)
3ErquSnF05CBzLAbYVgAMube5I1MpwqqXq0zXeXUoSDJJMkg7c41WODxMNddryhT
/zwEiunuxqkzM3rM85o4kVKVkML8rVdGMeDoXF2GmeLlwZX25SOlJud3Y4pRHbg7
VusJCflMbGqf6ab5+xCm3GQEy8H41SQ00N1hUNvgu82WhexqiazTSj1uDZ5gPEZ3
Kx3+UdEF8SQyImNFqi6xAejzCXSU6BSUkJ8qM8WnfLI8wHE1GpdMowBphA2Q6OPl
2VkNG+sefjVUOsoce5/SjBOXswQekZ+vvaVaA60Zm5/VQjjDejdRc0+pLq4aOhuw
MQ3D5O5Nw4su27A+g+vreTAd/Zk/RYuyGGiCwzmIednt+5UaFtbEp8xjGeKTZYgT
la4ePNmvsHFaRTZVXl7aoQca42ABFtebVaC32r0Ux06sGsxNhvHuVwN7kFPS2QOy
YJ6oPZLX/uuWW+pVJ/0ANwUuk+Q2MDYqUymZKWZBLd9xDp+4QaBUj2PZ17n6hxYu
nkbO1Xzbs64B+ZM4Tlc2VQe04S1gmtA5TSGqZIJ+cGLTcVhOLlrIMuaui6n+jhTH
wFG0/XcL4eNwS7unF69afFjIEfX1OP2rLfsUjhvTAX15eLICK63x9WO74w6rh2z5
1nR9y2qYp6QgH7Zve3a6tUo9AKekKV24+NMur2fSeiJNrRVNYS29mtZ7Hu86l220
mDUIhCsW8IB50w1qdW/aDQnnlVgectHqny+UF5bGkeQYTcAxL6Jsj9S0ahB0jJo9
tX20onSVj5gmlnyK3Fmon0WHqwmH4EhQ/b5bqDYuUyEMrfUazf+H1YXw+xDitAz0
Ixgrm083MW8DOUeyQwDmWHw9Jor+HT6gy480Pmo6tsqVg6aNndL48uyD5FpieyBr
ntgNZqix4r5c5K192hAZxZ4c++8dVL/SNbjJjzJmvMx25QL7EPt/RQtELmXG1D9P
GMLi6lLtVox+hsv8ToLmsPSa8m3Ev+T6Q0aqqcMT7cnrZb4M6C67E+mXYcKSg74U
8uKSH5D5F44s+vPFXKG9vGZgYt9IIj44/oXp96p0nEK4fN4tk2o7XfSP5OwWb0Rq
O7nlHLG2zBNlAwlBuQeusMiiI9cx/KQw9c82if1vaGOT9LoAGW6Haa833fSA0i5i
EsTdDujlNrAsoJQ4GZOQZ3/bSCFfA+LmrfSVWw9nDJ7m1rLm1U8V1wrjq4ErO2rc
lWHZh+NwawnP1U9G8CPnDRzAV4p1kykBb61stxuBmaKMzG6lrvWuI2pcDDck6K9R
m2kbEk8SJNw7Hxwx8FwHREo0WYAgflB49F2fZc9QY+6fos58+vrznyNgphQxOCOx
+rCyBlW210QJMY8zwRUkezw7zQv2Awv73piQRkiMgOqkF5yG1ufL6q/+8LhH9Wtf
vRS3zkJxVF9BzNwf6M5Xx7hwQuLuoEywETukMVAPfhlknHrhyGhdrLCYWdVDrjTp
6rH0s6+M6YGeVP86JEo/Q+/PPymNDHjxE4BSwu5JwxH2wp9kLlaycOrtFHR/MMs5
FrT6PX/t4+WL9fTcNMnNbxSzw97TLYdJxoEhtTqNXF9XDqcese9QOCgLhVgH8UCZ
2QiiY0dKIeEjQ9EL6LRwX9Job+SsoWDKxk2IlZEMm7Z0EGMBXF82Mq8gNLxv1z0a
XicioQ8XMvQMWdy++0b+CaDuT6EMqBnGC2hBPrx6Ux79fVsFDEcyLvZfn6IWAnyW
VUUaVEmsDYHIgaRWcb8k5CKNu+df/7btohjwUsFUS92HBd+blhEDNAiMzFVUsO29
q36pNWUMWxgPCk1RI8FCdu+LxJmjokAJFkoWWFmAlOMRRqeTsCTtCJHXnTVlu+f0
1fC45wSeTn1y1Ab0hZzdVQHd0fE/OvvRDff+aqMTX5qnA0zp4jeJjierymVh0TQQ
CWpghIMUcKjB0rUvX7Te7AWw5EBOFKV6y7JupRo85rXioD29mUFkiARLR24NsaQb
tTbQoJcrfZW6hXw5R1Ryx/b5/zg7x8Nih/txNdizyEM4hrpY1U5Zwbl+obfCSb/H
6AhIQRX3xRkVWvfa0KB90ERbxyITyMhEy8wyjIukCu60wGjMmzpoynps54yjj0ru
iToJc1I9F0bUyB3fMQxScfAlAFw65IBVKM3iLPRq+SmYnyEhuu+dMJtzskDWbPOA
7bvkmDyzkfFvntULWfrxTuTUjJAQeZbtTKbWLU4ubvrzVR/JdrgsbBPDtfh3516v
Vx6N7kCAlQue+eA6vz2lNQR1wgVGHfRYlsk3kBiiZsxVO4Rmm2oOF/pquSim+esH
HDR5yx0VfXO6i7ZAcaACkoEf9cDd8RrPD/TV7AYrV3iQMmoqf+lXMvPvn8ID4C9t
d+J0/Xv+3rUN9mQ84g76rbfDrI5Q8Cz4ulK9wT/K3366SYm9Mh6qgqR7+YDXpw/H
Mrd6DVaj/cyfCs50p9MGUmNcwQNVEDVfUvaDOgkt291DfjHpZCUkLH+ylCmrElAb
oCCerKYLcDvu7P7GSY0ap9jUq96U4I9/dN7mcaRfvzta6RSKykuN0LN0tYJ2lu/i
4K0Bau6V6N/TIWN7HjhpfI0eZxz+S/iR7FJ47619jubArvh+YK9974+v8mFtSa5n
8k4xCRintCGQGTLKVx9xEUW9awKHS9YOOS5Ucr7tLDfWKHFTWHeQI43wY5w4w//5
2FG+xxpqeYBqJlwG+zltYdNeNheYkfk/sQXaztht6J5Dxr+uFs9Nj5LhkzbHMH3I
xCFSY5RF+aIkmW0vXg3cnzdVOfOU5PriDB0LBaykI1JMCkx/90WkONqvSe2/xIqp
N2ZJYT6RapEly6GB/Hg10fz3Wpe9M6iJ79WTfzcFXbSh09uMnPTRzE8KvCqByKD4
/aadwznJbBenKlmpKWitxrxErYaMZYD1jWCOKQNvRRhgT6+kudrn5uDBEOCI49Tj
zHK0P9het5CLwnPoj/gisBJQsTCfhxY6s2nyDPWMKX4QQmQgYanVsbqmF7UPyYs7
sCMIAgaKNxCY91uCKayEoi8i8TsF5WTStzgT3inXR7qvH8uaCI3A5QU231g4/W51
t8gwl+FX8MTqOa/o8YoMuikwDm7kn2KPyTnr+YGJHgO6cMmIPA9ga8nW/4kIbrXV
in+Rb6tvvGNsS4LU8ayQ8kca88OF/dq8IgRGno1cxYQ5b2bOTo/DBW1WAq9mt5OI
p0Xx2pO4fDpJKmXh+/G8bdUy5JylXXJblWSRYvTs2GVlPmCDY6S6AdLnWCa8XOyP
2AkKDeRmNiLyVOdqkn4IMJMgTEgHtMMXScoIejQsTdSHVtZMSZjwhL4goFxKBQAl
uZkzlMLQk3P6BzQtAmma6gW6bxOu6ofnd7gS/ZUPY1M3y44ZGm0sYrYcTiJeTOM9
yshjMPjIdq9XdmwA+bzgRgqagkOx1r+dVCt2MPh97lBjcjFkOR2VCEKb2lgutSBD
9dT+wSfAx6ESZaG7X+E1QK6eOidD8o6OzoGD2F2ltYzg/bHOtPz1xGroSowbj8Ox
p1ZKHd6Zl638r0s57RLF8S5NpLcigCWCJKWNILF7WdLPZno4EbTdFj9Pb6usyxwH
eF+G/TK+L8fRtn22bIKQUniGQuKeTqlypJUv7VXyAvwQd3qa075eDLrWzN/cwNG/
CUaKpDTOMwrKYrJ68zG2nZaxTXwo9SsxS6j+onLvZYwPLbHhEdJB6W0obnzWYt0F
c96w60yrZlCjkWp+Lfl1ypvK7y32NjoavN89yX6ilByu6FK9wrt4f2TsvKaJLduC
56LYzSp5oAsTI1nHvkOWfAnlpy5e6UXjQGPhtoYDvqKU2D0iFQ2MD/JtgUzJY1gS
TDGka3K+kpObeDHFBu3qjjY43oAAhNccby+Tai4w0hPirUnJYDqe85fWHSIsDvse
zy738t+T/mCg3ohy9k/J1WhMhwr1nDFzKWj0f502JV1++bVlskLFjkzMXxJk4NJR
nryn/XQJd7qY+vcaOJelSohDVhx48lL7BF1yvBUP9zA4UByHNpsT5zvEWAUN7qsL
FgAnJQRJ2KckpiV/rNEo9eIlvWan9S3/n549Fxyp1bwpMDLVABk85oGO8wOSsz7h
es467oYi+Sp+bx3h0YfIdkGmI3u43wAMJ0lBWgcrdrPlwCqkV59eI1riYkiHx6PV
9kaXC9eLfx9Kkg8yIqtos0rCaH0arp0n1jLgdCVaKCwVpUQiUca49oBDWLTrdRCZ
r3jzSdGLoaJr/TF6XNQrqd1Qz+rXMOgnPVLb+EpwQ3qifs2nAKC6CP8dg4K/5cyQ
+9laNAtbK/mIeKRVWbTUGdlq5CDlSuhPZYeHEhd1Pkmet1yIi6hBV0/IV0mp8AdN
JQaEMKZkwRtgix3tvq0BGHhGb23HAXXWDfAWI9JwYS2UgBCZ+zDmjteMUBs4zNKH
WZRiFeJQh5pvjDqf0M/749O7Hie2KAA+rfBc8wTGuhz+fDQFBHWYxNY5ppQI9o5u
hrnNQCyngJDRYk3vBM0LfBWg3JA5GrtnxHRUer+fk5X2N9yc8tjxu86DeK0NoBIA
6L96XPv880HN5Gm2EAtCA7VgcnJt+tNJqySpvGl+fLNUqNrlBZape6Xn7CEqfiBA
592VaBCLGBBXPv0ivtuRX4zy3I3w68zjxOx3Sz86LPEB3aOfFK4u+UYyfSv1iE/r
3Cd/AdG9XVmHIPdh2+dU/OnQh/QpHdVUZJlkAk+07gf+p38Z/gl9uu35i+TVYe4g
7i22NPbdIDSN1idIHFwzaue55veAV/YPcv2XzrRoH0xbaiKyPECDL/Q4aDo3gtOF
TPogETkrovZgKN3XJw/v8aVkXdhucVXJQmWufe1vbSNJOGdrZXyghD5GR7S/38V2
GKHxAcABvY5dGHe72niUoaAAtMDmWZSuva+SzydoyrMMWldV8XEc321SobQcSjSG
r4/s0XcY6a5FUDa6uFoRBvMsrMWs8/lew+TFJXHYv3oh7QjTn1QG31Bk4xdzphpR
Zg6LvasQCbQPoahKyeURZ5TW3CL8F4NszeYp6WB3nHTjaCUyMzt+YoSGbgGn12ZA
dII6FxmOvnYyoMzlYeBqkvZMw4kZpLa979rlBVGYdTNBZvseWw/6MarRsEY6wm7S
6X0ddQa3tn9glQ7KtmD5+jh33Uoyb0uMEJSKn7AGMLWOqUEu4euNAAt429GScGw6
W8uCwvGKsOGfnXYsVgsJ1a4VhHoorwd6s7y5xJ03m1Yivte7R94/8irS5cqbfyxU
2eDGmcFaBag+tXhxb8DYJ2WKDNtOWdEsxRJAMCttFlXz8CJ7dG9lEpER4ZVniBWk
sX8ODvVbLtvBKaYxDsASni+RTdVypcK65H5fHPBTKIKoXR8aLs7HpD83Pyfp4BcZ
hlHx27B5vTd2ti89A7fEDi327k/Ouwyd7D8fVTv7UG664dVrL4nIkJSaHaKA0w45
Qamq55FcUVwqJad5PZ0utli+NH+tv0H285jr6+kdkYF2rIdPsjePL6ai1rKVkuaq
z8s3Q9TrXlSPei2+/iNUexGcTXA4V2koBTSFiib89BvrlgAjcN3EsCdgwMtNAqsF
7ffrI0N4clgYQ100kuCJtkZVmVbPdpGlqIKa/ylba+Uqm+bzllusPjwjJOb44zvg
N8V/02N/d8MATR6HuPLhLK+AzSOpBugf4Z+s6nfmhV2VCUDbWhqPk5hwFARTYWhY
HXbmame6fhYBdO7UtThbL7g9pKXKoLEE5ypKs2czuPt7GgUevT+9kmzJAPL/YTUi
NdUEjaU0CgsXVfX0w1B4aGyaLIXUodpiTOMfD+P7ohT/G0H68z149+4icAPfuaQ/
8Z6vkIxQJ36Ao4pE99kpFtH7JTUOEvl8gjpU4s43APGBemC3uQ5wbjSxeOQlo1BT
INXOWqMGxol1tPfSuKX0qh54XMOWGzN4OLX3UbA39hxW1JXvonj6reWCWoAjxC2U
YhCN/a8Cfp6yAPKs8aDvWMB5FSL82CrgaYwEM/7jVlswP7gdW+s0idE3jY4Sdw/b
EORwo68xmagwY0x2zXPNErr0X4R0TRMKZLMKwxqtkznf+DrD9PN2yoCLjJpn+kb4
Ipe4dshSWE2LiKfJ+uw9g3TgFS10tyRQ67ylrHG2EhX0r7Qb3A4VTlRgZ2b03Qlk
eBLdcE05WUwgY0j86ocfCLjGr+i7uwcczW9XTx4h3lzNW0PCRbn5QeqjEnUP4F8M
5bBuTo32YCOlojRfzs/w5U+KcgZmoDNZNNKfJs9ufU/7x2Bm18QVCt8G37JTPrph
FI7T91W914/xYyUKLP1C4nzvZHSgxc/ilPG5K3GOUG594Rt8AP8U5UVVLv7c/Nea
YJ8gkK7r+yiitFr6nLWgvJzw5lbNk8lIsUIQCTzEjEj90ppaBOlhtk//ClhpC+Ud
/9WYQ2C/XDdkY9KOI9GC0qgteJoDFKixpcvfryquQryMGXNenNuKrEopKSp56sNd
eOx8Eqd0eaSm5qvYLfDd+yf9JFFulbZ9lwXxW/IlpRosPp5iSdtF39tUlAl1d19Z
pEeImdGmFoZrzARiOey6NQvW3KTC4tw4QvFNP5Xxkm+uoeAebTBH8S64PXfeyqDF
r07AEUPe0gjTARwQ7oWXzIP9nFSToowoDOzqApn0c/0A41ZFyY1+aqBqtH6EGkEp
Qyid0H3SZad29bIWw8PIO3cZuUtV0HLlXs9HIaSufiT9qmU8zzt76Cg0CbVZcCdS
cvN8yRZpmZ/ilYtTb/OQl0rzyAvsyt3ZB7UzfkBkW8zAmcpsk/pHb710nslqMFOz
SZwLGUr5s7H2OrECV4rJWMq2Nfhk9/pOc1ktflSOOiNgLEW6fqIpuUeN/szgkBrr
FNy5UUC6HqDJf5k+42sKn5/8M8qkVbZh0+un00ShCiRiBdmIA9WCnybj5LgKsT7c
NpqYafD9HQQjlbRBoXPuXm6KOvurRWRaw6I4KLQwLlWK0USthKos5+ydUM5fq0MT
EZTwU07d0u7AxV6LcGhSX685bWSaOTvtidsXhdE+yXT5woJeuP2Q9hTfLppsspJV
+NJwhRTP3H/sbbAFImOXETA4XuD3kq6f0vPNfVgIu1ZexVEGMACiSlXOJ76PDMa0
gAVaN1XqcC9K+Jf3RFzYkkCUqc+9QTtoFBgyx+eiF4aqr9iFN1axmJCCQ+c+cetc
/xX1EslS0yoEL6WW4h5+DmcfBbXyRaAyGcyKLOVGANyELq4Pt5cpdXTONyOUuQpR
WIbN6FoHCWQ3kKTMAydYxUcGfz1VkQtT8hAkjCGZ4PF8OX5twaxPfDW6OQRszHaz
U492rqfXOUJju/xaeqQOqnPbbd3kG8ID8dJrfoE4piyMvlqtlEEX/5cmue+DqNqI
AYvIr9OiulWyFG0UzLsN64irI+TNvbcefpmrtgDS1CePEjex8y98ZbdRhA4z9Bgw
SxZEi4rTXgR4/TpMYMLdvw9HhCVgYUC+4W4xbbMNRqWAzazAck9559UXLC/RKYWy
He8Js8XSSTr6V4uUd9YMTMu47xSklfYv63YTCROHOkjYHlYvknAnVKDCoIakFgde
Y6SfTmm/BJImSEy4XyAx67tBai3pb+zSXjJ/W6/1tHLsiyaxNwqbdtjDvsqOZbKC
9KonoY77pSrunfG5EyWNEEKz0u/MI6DY16HoRM1xFFAtxeNnHKnu/f9gDn+a22Ri
JQEcxeGvBPxKCvZTrDp1HfcbwEHUt34hUt7rmrl86w4GW4h5T1o3hMbxUQ4QcxUk
SjuntSncwJwVY07sDHmdQvRZeyCR/jBk3VfDjrp2HD5qIercTE29jTbJP+GCtawT
DD22lYZUXh38fuZ7b/+2cOKeNhWG8k/3cLmjnF259xLSgwzV6V4VPIpPKCD3XoRW
zPim5rBKwbElD4vNMX833vhXYD0Tkxaa9PTvUboTU0J4AYGf4BDUPsxGnPckAsYS
4YQiAy91YK9NvrMVB7JgSYLTbnGJV9s5YgczfoVIMTT65fI40f72KauuYUHrMNc/
rNOGrVN9sKm72QU5wAc0Y+hI0YKJC8EkfE33YGdRWeHvEO1M7CUPJd1R0JIt4TwG
xPK1pwig1tD3kCVO/XEdC4hIVMIj1n94K91W9xQg+XAERr7ypsWBhmKgSK7duf2G
H51DTjRSxfR89D5fE+rjeXZVVSB3Lixlm1DVscuBkPy0L0ixSL4jDlyHJl+t/Bs8
s7bQJn8tM+j93r9/HI/uCrRpaOjvjPH2KFcsJDC57RHKcm04FKWI5eo72qDY1FuA
kHcsuHSprcXiBYbDx2L6Q64EBquiVWjkx3vylnfWir0//uP0qv/Faz3l8wB6dt3S
nfhdvDX2qInYp9mspKXzOB7TIEQMvhekbfzV1jn8oEcHWzOES45oljRfp4syF28/
qOCwhpa3bdOdGa3TOrSmJK3UWmbLYb57Y9Ys9HC5rheYNsQtzDq/Ss3WsBgAbQG0
FsPwcjy6XYxHbQy5OzifrXmUUufLt3siTmC6NhpoUwWBr5unwGztJ25jWCK9uktJ
wOGYX306/sTBdm3ts/ARXc4CPffJrwDghPJ0Mg4WfNSPMeyYf1BAEo4r+sBUX+9d
CPoh3Pw+sYEL/MwgqxZXG9ZpnswhAKqSettCTqwmvsT0MJlWY0FIZQ60mOjDWfUP
7+h+GVCgoq+DzQcFIpm//Le9O3+rwSsZx7fMXpkKP9Uj/0XgJFtNQinBN1H9vl4J
jG1p5uPFJ46GPvvgFciXYZF49/CgJnVUp/ktcZyRvP5nxjFgtbKK59wTFtCQCDye
lgQyy8+Ndv82224UYjEUxni3/rdf3YIItqg7U3j1ZPhS9QSVC5wnl0wJJLtVwRTf
Po4XXSp3hpweRRPVyIbUHH85A59yrL1MbKsWNk8xxinqsoVIHnq+ufrtSdw4Un1x
P4tHWZ3RIvQdPumYw0vZbVVZIwgrj3sTCrPykLaAB4zv0zxRK5VGTyKrXt1f2+/z
Vk6dBbrVvRzn/bvQvnTRC8h7HuPHBShXrXtYJZhTl2lHOfXncVR1Daqv9pOHvxCy
NCKYlq4ZX3sqY1pNPEqQV/uXhX5jEm0LxFvjKo2p4Ibm9bWveI84nBuPKiGAK8ra
v+VSBKRb8LnxYu8i/KdNuUEdi7L2cDAJ0m3fl4g2Z94yuosO0ooY0vfhMVacVJxV
9fx/F+qzPnr7qXmi0DsUsrNJl3r/WXDWxC7UCcz0OUzC1uAlaZwF4ieX10mJWSj2
ONqT+GH/oZBDnYy3FUkMTQ7r+Aq+FJgjTj23bFK+54Jo3ie6SNJ1WA0p2bRt2Oa2
Lcq+unfLoMobW40xRW6ruEiDh1eRDRf+jjLDqrdMvWDKK4wZ+eoct8FELccr7BXp
wOynwN7xfrpBn+E5EVU9qxpKsqdvWaKwX4EhfVIQOGiB2JNXs9DKyPGWs6Mad+N1
f58atuqmJsCTFV5/qNPus+n85z5xETyRAkunfyzlKU9NAgn/HwKD6UQHBxvMbbTi
eUu2zuWs99xqyZ49uFCG1RSN+Sve+yhvk92gPc7qGbVnvjzEKm07sOS+H5ehipDS
IbqGaPGlcj7aEn9avnEc1y5+fZcpYElZcDyc51wWbvao0dlitshu+Cr8MguDORKl
RFpaiBMfnHLo8pPYrB6Duu5rDzNzDH8gJlEOi7COu88GoCDwNpN2txw2+ZJdZ9Hp
mqANTcdMbJHhB3MkoFTcryK67+gRm1kZs2yhaQ0UOMlof3xDanodBJxSVZdZQ3Gp
kAXgetg36Z6N7hLLR6UXEOHs6EntehC1L05Z/KTnKB/Z4sBkyoINCPDiijIZCuaH
v1RJkRbfvbluEWcv7iUXv4A5Q05pzguoMcn3AP2kJ17XrswQG5wosQaH7bNTwuR/
k7H2gYxlS/97Bv5RNTpxJe1c9wJ/vlSTBo73XSS5hOjPel1ktL+Zz/KdmCfngWGK
3w6KKPL0bc92e47hh1eYElqI9dwYXPJDKGySjJij7iN/YUYGUrQE1RlhfyCOVhgZ
hxtZ5UfZwHdnu8599SJLJKmVMBtFIDOjKZg7PigL8swDTJrNCwxshcLEoCKJakic
biU1yl6w781Rsd+XE20JUVoTH9jT4/UwbN05FwGK625G7lmwNm8c0bDQTJi4oONp
65V67jInmN0S2u/ihZmTDeyVrkztnyQfcMWdPFP3lMW5xzUJL7mJ9gghsEovb6mi
HGIpodQtYeD4+ekWf60QOtaboZ5KFksAi2saeve/41HkiFPRv280JDN+asAXc3Dy
5CZL24IxYg+HXn9FT+l+gld2rNnFk7QxnygMMjFks8dxxVUxBfnAkW4RzOE6ec8N
R/uxmvXpY4fZa6TKx9GxmsvjmPgfIchYwbzou0sfiEwXeLGPxBeZ9oGIg5Pq+dpo
zxgmeeyrOytDXAi/6w9MVNYQFS69PWmxrn5Yms9w7Hcfj2kUFBMABmngocZ8mtHm
hYY6JeK1eY94aukvBXarENWAh0ZdtOaK6ykz4IPKw0BXY1VsZrXpp3sTA86HMdMx
bFsoxc66gzAoC6VPgK1lwmI4XJlW6FLYwXUJUhKQtJMhbBfWOiVJHxTOxWXu+deB
oH9jkYLa4KMLir+87o1Sj5kmvZgD0ekvXgz48248EZw8zWkw1CF3nDaOMePSUU96
SiYzPGZWHXu3KOGJBfmSbIiScFJ3kqIHC2DiGwaOrRcrG8Xp4LryWVH8CpeKCypA
AaJUnsFt/jAsYKuhm4UzO7q3384L5Ff2ihAPjy7imqT7e42XSyVuNBiX51D43qYn
pVriCzc08BD6Z28gsLT3yPosQKYs8AdkEcA9OO+72qZqEr2X42e7GE1oWzrh6oig
DxC3znmOYwDxhLq2cg/QoFyl/rvxHWKgUvsjVp1qBnHEebq4gqpD8vpjZwrvY5Ta
K6n9o/PMnouW5fxrE+KSv8y0FfrTTMuvLi1yduomwmIp9FsVXejITO4BI+okIsdd
wwRtoRjIZ5R1FKEB4Aim038zs58xZjwomJF5LeYMeMAGpiBnx8LvzjNBBr+SvsYy
lQeiZfuGWAEnryRxRFqU9cTHlXL9OGy5lqk0d6kDLWzpxFrxJ1SoPCIUfDtZQm1W
pv7Yta1OtLAQhg3fudgl4yLFtJoo7DLaJgbvgeEqQ5t8USlkGM/k4VxsdXEfecni
grHxRRih90A8LYmrvioKPn2afAiR6MQ2uAa2zqkZcBorSWpueGj8XDlQ6vKElu/m
w6jDc++CxogRINFq1HxDrAvjJqBCcwdkB0Nrfuql2TF0Q3pYPdJIb9ZsOoOGNMtX
vylyuKsiikMHc/89KciwC+dgcJZ1cS548+GDTXG4p5/lcYBlk+f5B0Sc6sAFPwrX
nRpqYFNFGuQ7IV3udG07L4+xRBwgPND6VTzyhCiJeutXUPDF4wAAnAPZ9jFOmOsh
UoHXzpq6WOQoufiGyp5FevDmkz69lAxYJVv+N55mB+rqxSfR83cYFBvuPVaeSa/B
HJuO4JFabrCsbDSKxv+7OLsYkZTKFsa67xxj/zyAadDwmjQsoJJvQ2b1pTQ10ia5
xsE1wGBkqBftjJwwOXFrbHSy7pL6nDM494OmF0/TpCu/SS+eelwvQuw6HaxRbkOP
j5nXqh8lwhHg1DoYzVItOIwqzZrCCSWO1vXNoqmy7yeAWAf0Ru3MftagXTyzJwhU
atAh9WhIofPsCAPA1BMaTZUAbXweRS7firAEa1FGaQlxWvXzdKqlVOXPU1C/E85l
cn2+g5CIq+HrcmMPBd5xs2sjlmaD641pERbt/HA4t6mJ6XsrRVL9vRIQQyX4vy57
FtJs62WszsuOqVvauqlhIevxcs5wkMZahIvjIn5i8lbHKtfDyTsSPvy5znfLbcdL
Q8muPRk3PSlR+jiG4sp6pZvuEEiZZXvGjnVRTmalDsO6/KxX3sn9vfA4XMZgY9zV
IN+jEEPUVGVShCHExU8ccmtEMOt/lR+e1ST51Bjfo0IZVBeBjBcCMvKbPXTQaW+8
L5w7H90TTJrhMvqfOyoepv1vkjo6pekDRUXFvQr73JWse3HvxGZrLRf5aNv9enJZ
WDRuHthJx3AU/caTIApc91367Qn9IZzzD4XIh+2EojksOXdCyZ/uZ4fgQNUyE33H
d37Y2tapi2uNPVEnYErHjVsnWPaSv1vP1RVR2s/aldfjdVssyA/v0wHDe//VsAW4
ukF+Ctru+Nf7Nf41DiRB4Ny75ONC3LlNeQ4dv+ky1VZ0X9jLGB2iXV9mdmP1ehwk
ruiB4Vz0dg+EbY5iUW68Oq2Zr78sLlpfRlGYXpjVcwidlYb14+1eBdEYn9YKmynE
SaFBprET3tew1g3x5RD55bP+oZbbqdbFGkM/HlirRYXsTgcXfQPraEzj67x7rQf0
ETVkF3lBWKt71/g6ZBrH4vgu5EwetIwBkU8gIl49Ms62WFUpVqRGst06Yu7FHw/H
N8wAVhkytQzASss3y1Dw+f+nq6wSaKiW3WWPbzGrZ49b5pZl+mVqUwEDGDufV180
ja3TaM7t1E0UhRVuhGCY/kZGxDtIF815fC/t6AwW+eN+RdPzy3wNW2YE7i/imGnc
DTqe9gfHNTVEQrEJ+v0ILCO458jnjZr0fEJjKu9VV+XB2LpS8qoBbkEQI8w9Xt1R
mDQGb/nW6GqeQuUtU3fW7Yl2z7qeI/geTLEUukTsPD9ISTa2zxab6SpR/S8NNvdx
+t3pab2iDhxlDWVmIBtM+xzsi1xxyYfQ2LqjPuW34rEXKGD1Ynj7hRt1ZzX7bX+V
3Ii2GzBAnMs4xGKYzYxQ5vu0NB1zD+2Oi2PoyfyzGLW55SNqUlUW08TnSQkmKXhr
89zBhfB+hPzjk0T6XilPzDprnMSo9omNY4XovMkHmi4R+VHJJjqiTBg5B/MmJk0S
NPcnHDyYoh9KISy6o1Y7mIQ80JqMI0mYT4ayFS5GIRj7eZgZ6Wz+Wcp0RuamQLAH
Zjz4YCCUd2u5aveHgb8hWv1N7IBF4xZx/SQpbciz6wA7ZX2v1/4ZeyuFI0e8UQMY
UIi5MN2dpCIAbeXSo58fmmFKhD4ixyNdNsYdugROK1biKtNjE9c47tS3Z2/jfypb
CGBbNKtRQRVyU8w8W3R/gIY5sMRIBaErfzQShIKfyrnqmmkjO79bAOd8IIdmfQ6F
OYL6qycSHcPClafF7yiz748j1/7e/iCerpktU86laZUN0Vryn6LxsNdLHUzl6b9j
Wj659H54T/5OLXfhuQ3DKpGgHsO8fuC9b+3b2TNrROAIZ6Xf9w347PFo6/Srhnwm
Ifs4sOUOCgmEjK9atrY+N/qjiyyEaqKXJx3V9jP6qpIU8sMoYRbIK5qgpk9qN2fw
ZcbB8LsXLKfDhOoi1CtTOs1VNhqkPQBAZwPnosT1nWsF5LpD1tDJxlp3n2y3hZFc
cy2IgyPqA1oebFJB7VNkfHRe7bmTEOnavEzplgfmhWRDl14thWHvFDeZNzQwwMoC
pL8SGVDJqDiF5CaE5xeEYMRWYc0zO8ecKticqVs+gP0JY83FV3EiYzg+l9FKnzv5
oIhThpoeK/Mf17eUP1HKsWn1VDps48bEKlNbuoWFrEluvI5VsbL+eUYASVWp2p8i
b/D38/0ztdKrkZYPX+gA3xN4+DyUuCxVIiUjkqIEBp5wv3NkaVs8V86xvdsVMF/G
HMETRZruKbKa3La6Y5SAsIJYiCsJTkM/9x+xEOFdMGJetE86UcGiFd8aRIMz91o0
/Ldsbk9r+kx1lM51vS+9urbJYWH+ouIHjU7ppXB4VZOCql3MuEQBiFw7FXuVS6QQ
7ggFu1q9w1hN9rD1cJpWaSe+jdrh5+YSNnJPLOCejDRgVfWP0taROOlFjYEKCxq/
DHMiexpGU54P6hKNmyGrwS03R/gj5lxpJHHY//sjgorexdplhVpjWaTNnnyYPwvw
Pi/9vzcAikaEf6s/BmDI8pWc3tthljAmtXBZ+i/D5HhhS9T2BTbxuB9uxLJsUmRT
Nvs82B9Qio5+Wh8xNkOqBFl9IBLayut59uKTn+Pifxo56rgzTCsOk4Vrd9sJMwA7
Ems8X7wXJAITpdSwNdbJ9YYYqGaJy4r+WaK+ecDl4OpPdXCzSem4Bvzppa+zH5I5
gIZ1ZvL8yaR13dAJGkAmA3ZDJgu0gkfuWBoOExZs2MnCs1/hNLIjRV1jHyhpvSgh
FcZtOt2UfBm1LTMa4CIYzqpIj6zLBdBV5FYNBbJqIRVX/OMTDUpgAVCPzL8iB+OJ
J9H31uRZKFPP6sVrzDk4x32IrP2pCUno4Zq85l9msB57ZQy31vG5qmsEZSE9ljna
mWmFoK+XHUM1vaS5e9gPv9Tl1InrRsMfyJ5MfS7NlDaggaXCCjaoEHAq/IrHHEdg
HgsC6+UtK8UmXLgQI6ckmQr+gi3Lvvn6jTir5JFpBOez/RcCdsEIMhV2+ZC5SBMQ
umQD47l5u5vg42qYjlgxi4z19xLEwtfxDbGQVlYUGOOMcq3nQx1Y6VPupenruw3p
dIDY5ZcZyYliMoyUgox5QRLYhA8Tvxvr/HY/+U6NeDTBJWlV/i+qEju89Un2KEzN
tOKMigEvgi6EOU+KBktBBBY5dTYdk+ftoB45CJQ2NE7w41DtC/wgbOmuBRg9B8+t
hLY0kaAJybm7Y63Wyg7vJkGIzqKBaIpD/UeYqIKb8XI52PPw9Oo0Xnsw7B63C4Y6
Tz0sBJz8jCDmxDnusMmvM3iuFs1LkcxKVB6gDHieTxd3GrvaTvM76VZEM2S0Gzcx
orNeexi5wBDbucp1EMTNf6qWOHI7NYRV2Aqq1Zpugp33A4JnZ0b8pxPLIEnO6XJV
MkCrvPNuzKFDNY/AFxX54Joj4/ps9mWJ1p0+Y5pQPnD9a9MWVxeAa9WkNyDaxIsG
HusysTFQpaciFz+IW9A/jru8MVQfjnVRpiPHzuSOYMtIZjqwKumVVESwT45Ug1lu
EWBRTxPMhI2TYDpneCWlAFJldRa+L1qOlypeIchLzcvtAEGUwKjxGAaqO1QdRSIa
a9MwBKzqmc96idqFlKhfyTlm9KlU1sCfp+nRsHBKKArBaZZLSbmLkP3Gf69hUQ1J
IZU6fxcZCW94vibwjvePo5X8FEqAkzMO8BFQg6qeh8rZPDtqknKIRjkEJJiG+Ksm
eb/3RMzBj/fKu50HkhTnAK5k2DPExC4A8mXdClZVidHdvdWqBCP+wNtawPmgZGCA
5iQYL5jxXFA3c8SPsUw0kxuWQuowg7R02OmKPt+97LSVA4YbW9alT8oKdUCkymEq
gSD3fxwgJzIJ+6GLXJfZJ7kpA3JtBDXPAktu4chWMP2Gfsd6Iq1OFEp4MQ2nywam
QaHE9tBrz1qq7xenKgW1RTSra+EAxZoylfPqL/9gfvaJ71U3G9ZP7I8HL44hRWCw
XiPRU3VdDMUPD/Q5etyf90pjjlQhWexP4zaTH3ydrL+4WVuRYSNrIaLQaxgzJm0j
sqrbntC0dUdYtr0ytTpW2akxakFnksolByEyjMS95XHQ4kURtn6wZqvNJuJ06wBY
PdoF13thkFQ82A2H3wfYwTuqryzfTtH7GD9wTncGbaAqANvNBxsrvX+o3aVf5ABZ
af7ohxqjYWk+2q2pJrN2qnHXKsjdzdIHVculkmNlhPV9GAqbzOCdeQcWw/FR6wcI
NfZjF5KUDsOlLGb4xBkbq3k3rEStwwvTqo7upeGP26T7/3F3mp0D4AXgIkXqwHCR
yamudMyBe74n0kIZT1xV0Q3AmeI+sAvIRHXh20Eizc+EkpNFBUgXq/jPtocMbRr+
k/6BkH9+MfHjQwGEAArRdObLKRebXXRTjCy4mPFuuWsJ1wCLYjwXeki5Mh4liHhi
+iMQJBzNBrQfEISSdDiuYdTe8BGnFyjZSr4B+JdEMDazhR8G+pJDvStUGeFIW2lw
GA2WIdap1PXhCUD95jmzebS4wL3efXovQclIUugeAxPZSawUswBWTOoxwjjlERJb
OEBtZLw1Y4m0gUXzVtL4yq5uHlwShYaz5LF0Zqul6cl8NCyI/FneDVFwecM+8g12
59FPZpNluk3T9hiLJRZyUKO+pnrxV0LEU9InakzrMlXx4HAVVNy8LIhX7o3ohAn6
MvjCfgQl9Gn822hVSaPYscZmk/LQunYZSgcChSvJ9LIS/7MlhcfCK3Db+vGAGNFf
k8nkpOYgLmUet3YO8ZeG9F8DFFKGBd0Uxaqqb8Mdha+Ixe1qqj+R89iHyWFdLM3X
TzWVU3eEsIJJyn9cfGuWLAD5w7b9r8bxjKyHaShy/CsznpJULUq4adRmmyEvjyDH
UQfsfnyRekPQdU+17WrcXvJlmXq7fMlO1AFE+w2Du5yohoPw/nICMS4ySkfm2z8m
u3b55ygBb2dlQaJ6v4XTNkb/VjqrMlDl7iPrkVHJ2264bDL7XH7KMTzXu0bwDyaZ
QyN73btQ74zRLN1WaF9W1sfgfyOBv2+VNg69YKOuZmwHAxdaC4H4O6AVHjkEcmvN
FNg4/2IUKcDG39K/L9oYP//ufX7KSs7ZvnI3fZYR328uPUKqa6ZnNVLcfBZrQmCp
arNKeoQFD7dHz9153PTlezTM0TDDKCQElZ5he1h/Uo/mUfLnwmJRkRZH9euh1U5h
zb7+YMp4BaZnH/SgNWO8MVfUNC2Mdw3Qn+9QwRLCYSuFpQBHgSEZUGKGQOMapxDW
S+FmbtCrNLxcOWGzFdWOhk0KXbAUaSuNz6OvCwryU/sBqVRNSkcP+MytddyiMrHk
C2dHFwr88d6M8Vstq8aU4sjDrL76+xAFIFw0Y7L9BceFud4bV4GtFwFI7t+EOxNv
x8Wvoj44vHhB8fIsmka8q65oYFiXlHXf/dHxFhZ38NWzrSfd/NHPKYK7pZbSWJqL
2s+BTPn95DAqds/iSeFtK2RKWBgfT4im71u+g0K45UYXlDt1JWGSDBbTVZ/nqVar
dZUulFd0rP9ito7kiIRsArijscCmqc+XMd2ljVU4BVssrcfZxKqa+0CHRwBdt254
mxmqa8IwL2WnNJZBGhYL+LYsBNn/AUb0zwIYi44BgrR/BXTQGT93ozCT+AOXShOH
nF0NDperQyiEEQJKVpAKAf5YX5amWXpHs+6j4RuOrt51odEfa0ZDcNR4Dg3O6Vd6
CS3oHCZHycLVoStIGqQxJQjr+i8v/89i9+rH2/eMfbwCYdl3tE+HlV/+4AKmtjMT
nSN4yb9abcxeiFwFsZ+KIkxl4Cvn3plKF1OqKJBULKbU5ZYACpKROjzHX8qE6YtE
RQ4SgMs46ZYhOwcylXuOS7Jkuc6bPcDZrHycp3VZHhvC1f9VZLP6wKTyO42JkMvs
7TKmpgmeeAM9kdHng4ZvImFY+KT4TUAhMkpN3PhpH1ZcxG7234w9pwU/LOhgMqTk
0PWbItGlRNJZg570h19RY5Ytdi9h0BHdX4XCZDjhm8N3RI+rNQiKL4oS6cmQxFZx
eIPO0LLSiG+91v+iDcz7pg/5rsEAOt2FWtG5oSY0gciDji44d/WV8IjaMtXwISkg
zzW/hW5pfLw3X+kXPwVf3YnWOJv/P3bdNe9GP1lXlKDoyHME3sXKgzidNA7aXKuR
NvV+J03YpB6q75cY5DOKw6GTC4HoXdvbIAZF8/my/q84QI9+jGKmZErHAJ5qWhCB
EbiEr+3vUZnxi5ApERt5GNRYxFVyDxThGcsf17t9utGp94Qfwm/z/TAVLVhK/3Ly
RTfkyrF3vKUc1BPwKoCMTjkKptiQBsf0sO4OOry88yTJraFvR+EE8IIPSW8v2HWS
CmZI5xbTLJV9PvtlHOcA2HNy+wqn6Eusv5s9228rzwhBMUgzUsSmIt+5OIkPiSIp
JnpxQCDIN7kgnjXG6QnxvPQPFbn4m/nyzQQruBKbhGhh7f6htBJz9qcKCVwbrd8E
uRD2HmU6VMSulzffkvh7JnqrVl6sNaqxEmGnMmP42nXNaJZ9hAuCl7/JeXXgVp1Q
clSJHUvs7JGM0czl0f62RxR9GMRWSGjTk7kj3QFWMrtI+WM/uxEZVHnyArVChFtW
BgZ+taa6ZX9SZSesPZXvRNHKR9oBzaLXNwfKphTi7V3tGMYJVgsJNpaVVVDjb5yW
U6de1jFLOysYdW1CaPtCljtbwYW7gvj6JZAqdIb79ZiJUhTNfiCnNqGbKpHqYqgV
xTfJ9JAIw+YpAZVaFF2dd6PKWPwANQ8hehshqv5yCibS6Me+Jn15SgtdCDpiq0Vs
KK8ED1qtJ1L+uvriGlAQ9komrb2VoK6X1Cv7QtdqP7TlYoX1QueQXBAjkYjmy4Rs
ZKdRI54xhgCwIpMl7H/Vfv5CyTgPwB7dCpzWaiNcshshsfuo2iBLgFC34ACm118b
TtJqnn+gMUJfo8QuG14TlxXXcEiwZkuDrIEvP1wrHwvvGwTbd7ivtnCwOU2usyn2
pgmeNh2g2VKY4Tij25tAvuK9wd8dt+aJYICQtdSGnVJoPnQw0xfjwgW/OM5vXxa2
gGRn/GnqSZ/IbEo39S/2irI1r9ef1SkJn7dO5jBiFZLQOXnrBpP0Zza99ntuu+um
EsnZ1BgOccKbvWRuHIvo+GeSwOS0bjDbjyYrPXQh+DFjJAD6xa1Cb4GtQ0WKi8LC
q9weMRjimjIr+xEXDyYINdUcoOFm4VHB1GzU+cH5Vbe7nnc7TNiyAK+8wLdBnBiV
k9UVgfd/fD+b+JBXg0VUPAQI7ZH0VTsA2UYXzqXy1KEK55a8AGNzKS1am3U/butp
cTdiWVEjpsoU58GACSgFFjn6IUGaaPpwR8B7zJsVXRgCkSdnDJQkxLCcNnIwA19w
/vu4Yz++aiCEQ7IL/VxRSElFl+k+8RlZEjHEkznYGFyf5GlmV8R08hvZFuugaW5t
upxFfeBE+nnYeuPzRpvEBh0xRvY/VWSNE0gHLJKkxzbskX1nQ9k+4Bk0Oc7YnJgD
xGAZBSroDfJs07YryaMgF7Tqn5XYR6zSJ+kdzfKpU86q7qVGEra/5L3JstGmFGcs
1GAtR8Imj9f1rv0wkGvO39VBD9mCwBXcSrK+rIaz9a2K1i2kgh5loqyrxDsKzVmo
YpLe50iX7WBXzQz1qf2MH5vklDkmneX2JU57XRYvSPJjCsQ909fsX2pkXUSkqxnU
1GMjPRyvGAgX/DazB1IvYscT2BFJktEIZL4qQ+vo4VWX4iKzwowLJRtwFqZFwCcy
vdOzn1sscdSMJQgZrdRlfF4lceT+tl4vsYri1+gwwAONsx7NOqH1nc/zYQyZb5XL
vfhoKdy6XVCysvhhX9EKzVWLE9POylGI4AOuQXtk8/1UCltptD3fVwdLWZq2ydSe
sf9xXSiE+1vewaGYeV7wrbkUcBnl5JMoEL+cqL0TFmr43AZaahFzF7XD4ObS9t1e
+TUs3ZwMOkX2UHo4xapKXea26w3xIdLVgL1BAHARzlZYdToeETQcBrZFT9vXOjV3
MknHodiJ/1X3/agyoehPynfdv6Ift/nlj5goPyrCngg5MFtblGQp7hx4KW1/owzr
ba4Jjw/duBj2kwSZg2Oo4Polw49u06BYX59g7GJItmC5H/oLhWzz0fRQMwUdWbfo
zYP1KjBq/bbKOU0IKktL59VVDzqQUaAfIz4tJ7hO9DOb4yW41MKZ24QPR2m3focR
hPQiEFXn9xEGPQa4ykqnEXpkQ90i7+82VrsAzV0JSveBt3hO36Gtn5ncbSUaSxy1
/yUPxzXIKPgm4t/1GkkWO/IiIwr0iEkblubBLm1MRVcBGrQq02aBGRtNMlkkK/Lj
D+0OtOtG7MFOzkD06gy9mtNxAjjr/dfsPevYOa1wfPLVO9QHnVtNcGK+f7v2EZCJ
DEB5vEBkeSpZh6JuupBTSkJqI7nVCzbhAISE4/ZSBFDgF70YhBHdkRTFD10K48b0
OStYfTqf9IPhMOpFFsIWG1j+QqNVODnwp0MGNVNb+HHMweSPVaBMs2WDwKOauXED
RVBnZP2GUpokg7l4YkvsaNBS8IRZe8hsil72IJlajj6abgsAhwOhFoXjCqY8gWog
fuoVGDZaLd4rUBcTJcOkkgK6KYO8jTszmDy3KYxEmq5uDfSBU67wjBPPRpILRXds
z1xxX82Yez/5PmXHrS+V9iSLOVPK2Svy0urCvm7CRMHb1JzjLoqP2/yFa7f3A6+J
KPOMTMQAbgy20sa0K4ADRDd4owA7Gzd8yDYvC/R411JeHpo6KnqsPzjsGir9565N
/qF9IHNVeqPH9ARiuwr+2nhnr4NsNVQ4jirn/DE95XYSyFmrAwP/w9Vh9G4AjMPD
YOKoEX3/XuKEiCmUR0exSIcoVOgD4zsMX1dtv7R6rNC/S2FOFQH3vQsFadJVfGV9
Xe8xeZCr0GnElqzVPU4WvRlUjGKC4JPH2vyglCs4+b5o0NWwKuoOxqrkR5Z41LS2
KVv6HikKLVdOXGjFdI+K9dZeUPLdFawMjr5fvJhMskHOpzsv16iOctXse44vglQR
rCkIUtYxDKuKNUQXrel6OntWP1NxFk+bZbneNJtgycbWOfhEl1iJ/kf4gBQT8QJe
pMcVLAkZFSQqSA2SWSlevdIa17Wii+lzRYWDOOpVGGnPqxshp18BlpGnTzqTytEO
uucjKiR8OcFex454LimqslTJetU1IFPE/skUplvn97kKtzFWCMXRoZB8JdSQI8SY
VpiJEQV7YWeBDuNbt3sw3f9wihHO9FYNyh4Ju2uO5kiZbIdRGXqzbP40O0thHoVm
aq9/SQJggAiG19zgcdhonlRMXPrEDo7hLoVSQResoO+Pnzw1Pr61w0Ck9ht7Fn1M
iaRFE9bYGQNiq3LQYJOmReD4yYy+0H8Ew432D6zkK66rybEDhuhphDVQAxDw4uzi
eySc9I34OajWjVKXhN47dsNTny9NRtPX/JV6wZl5k0EuBTHIqFfAiDwp9ODMVJeQ
ElJvRpXgJIWaOAttpDwjur5niJDoGpaZkj8vR4QqJZ4Vtq+5CA4fT5Cyck7AP9XJ
DeWUg13LWAFCCq7Zj66iJvco4Upm/wMR2/1ZjqHR7680rM7tgcPMvt1MOvFVhdH4
78D5eMJu/6PMbiTbFTNGuYVxYbUh/3xdBOl19sTherwyrwqkGRCqAjCZ45d2iLD/
i5Yo91M13eweiHMpWbTwCZ1FMWJcrRVHecMSfMfP9rVUWAUaravHE7SbYkJqmzz4
DfBtBsB8Eq1N4ipS9gzrZqnet3yocMePi3HwG3V5CwPDWgQI6119R/7QsI/WmgXb
RkaicbOzvIbSZv2Dy0hn4seWbYkNuQtwFhGiEze24ijKhKR9KSrC/St9Blb+JV37
JtpXqg/qXS5Tl0kKzC/TFaoFwb2+663CWDaV7GU16JSWIOfnGxriJtIwuu9k9wxd
e90B1vX5SeupT01TaNcV0c4fiR1HWmcklsOn91LLZHfgOx4LiJEgQugb7ta0370o
5FSjtbJeXtFvoeuRin3Lx6Otd5CcSGtPl0jNX3fuuIjh4hNDpfcaxgNHSssfDQvi
0lPwZBDRk3BCf0Ga0LxK88I1SiMiITDyiG0g8Ug8LExPJI0zNELjBTEGz9i2dqs4
FB13mjlSr0DK82ASIkClYxNmZniq5ATHJ/2x07stASFuBsuHP/yALSu39iYj7UY9
6GHer84A6tooS3ufAn5dsRMr+fAmNNS/h1L5nGO4WLomF67bHrzDN+FcBL/R8z4s
TvH7MKF3m2EwvV8pKmWZE3IsvJyBBLn3SAQ3+qcDOZLLf+RWTF2D7MrveHy7Q1BY
1n0EhDyisx79uTqh1wAQ5+ppo9u8+TMXyZWfw+R4olOwnWoidggr0jTdGA+vh9la
AyhYBaAMNDUw1sucLpGxcz0bKFogOW+dLRc2Xo/YeZL4zLHr6GF6GYVYaRy/2m7z
UI20PkTVUMIJo8waNv60zb+JZhU2uOWQFx8LU2mRaFTIGko44KDDZeLwDYEZlnlS
5J1Q8pzWRDDaGYPBDov9f2KzJ2t31p7cmCvh3u+DbGgAd8qJPZErvwZKANkKnRZg
ZKt1GyDVwJn9H1AmCsRvcK1l4JlIN2Ly+pYwk6gzMGJmMKX0Cnk0mDqLrRUAUxwd
L4Py395q3H6SyAgEbnfYp+w9VM16eSRbpitisdl1ytkILzlmkiyukpfbikDqLlz5
gqcAdFMlYUZqfE81f742MpvdiSeJDvbvDFVfLGhjte/rAte+BB1hQlvkTCXXaJZD
LHjJ8yj6Nzf++WpNE6iWTtj9iowYetG/P/85n2qtLgerMi+cv2hUs6uOAeJSZXx9
XXZEQXcqkhODprWaSSOlmkMN8RgyOSnSd8eL66RJ39CXQY8Iup4tcGddrn2Sh80/
kjrRlehD1rbd4InZazEM3Ny/0kSzjwSZQbDP8DTEqDCJMIo4duYTr1D5Ww1AhCvi
hcFmuBdj2qrbgqXCUququ1a9HE4r5Nfnzpzt5x3lg0EYoIcpW+NH2gfSBnBqdngb
2ZUwYxkETkvFxecwEdbpvPv7QM2dAoXC0cZOa1+gWE5IgHnRiWF3FeOpfoZlPWoN
+s8y1/3+cfohEpqwiu7uSf8/aRbOD10NJ4YQQaslJvIToyJMoEgsH+sQGUik6n9/
cCtOI8Z2YERvVg8Nnga6elB20CRcZLCNAIb7/T8J5KpOiIRNW1Cuyg0HA9mgoTZX
syvAU4q2HLAWyebHerWzrNLLXKbfyi5zCX0PmT7k8FMIMLm8Nn+E2ReyvOMXUe+k
oWL132r1KWyCWEMx8Or85d50XmlH8DD2ActYWo1Y0FIjPtkxnGRi2V0BEXhI52Yp
tmXhUqz5jctmERK4YAs8MmJ/V0cHatYG8NbsCKwZDqkgNoHF/PS8ZJwjBoipsgQ6
Q31co1EmBOopss0CyWeCGyD7lIhaGzbSFPejJQibs+JSFn7C7w+iEO39L8jdE7iD
x6SHXdN9lcURTl5e+d8IFdH9F20hawJBekqETSBkrGq9YGnd3UvJcUNGP7bgAaRA
LoK3I+9iPWNf0P6YHlphJBsQJWDGRa2wzOY8V5gDnMg0B/8fmVNhi/Gn0xJNMCGi
oghNsQk334xgAvE5fMjRZs1lP8Y8cKkFfgJsdTUz55VnZh6iCoqDwltkD8QXyX9f
/w3xhOzgE60iXNKy1JG4hVIZySz3y6EweqJZcdwa4Rg/Tqj6m7qh+w5wFl+BvZAB
1QqHn6rIO6Mg9XdQGzmqCcYHNMRyGljBqSZFTQqDgG209xs+cpLCXmj8m0gyJbkz
OrQ1NFBp4RZWkmWFMl29lKKa+QDZ5Bs1npJoeLSj/Wzxpa9vSG7d+mpmQ5VfmF1O
JEcCYeVUkT99CSdM/ULfDtgYKY5/cqJa8VftsAHD4l84Q2GXFyKEc12nQxPigex3
hMo+LNFyP9AO7TORq7gWx4pIII5CweO2aDzEIODHiOFTjSdFyqN79eBSeLeZju0e
DWdWathJ0bMG1PacxIwOxc+bAenekMGzqL+cU2svoyIVvXfDVLww9D2h1BX7wVAz
fn9cJVPf8lnhj4Fl/+wieLtVd8fXtmLCHDXBxdrGKZ6AKqEyQTBkJrbiH+iPS4uW
F8aKpnJHxp1bC+flI3qLZtple37Cg0eDZJa0XFTQ7bc1WBLU3aq8KDYwZxiWYM3U
nuOM5iZ94Akp3WtDfLTkwi9qUkPo/2FadN+f61Wkv7i0xBC5zgZpOBc1dm0kUITx
utyYmLx8xRLBsubKicrWJ0Erg3wCMydwXxPrs0P+QZQZfcvdBhJRejBWiPbPNFdH
Aem7gmME5oQ56whetgQgUCZK1S+mE8E5k+q+IoxoPOGCkD7qsRFqDDb6uWhwJ1Np
z2M/urg0/9gN57ZFuwMQhbc5x7QVcFS8Wy+Afaa3gAATkeD8+8B0CZCItDNcZPHj
mPlrM8pQ3LM4s/DJ2I9mavQwJQhC4UuodL25k+YDH2iZiRHmSGwmvozSrzuOnSE9
RYNppodanHoCGCvRfySn4IU65vzXT35vXohvACwi+mKQeCSf8uJBwtOO95Mr/RI1
dTzYDrOiH77Y1ObBalW6NI6HZg1n2JGsSZyctPbzQTQrw86ovOcXk8cqFFZ4KlR7
nCvwvsW3PXz8oqbcwlpb5foEfYM83jdZVdIGlhROHu6gsGy2Q5jaKRLj421RYxOA
xtNaV/gXNCdju4IgRVt/UbEgrtj8hGxDRI6tOJGZE4pP2zrPiNdCQbZAKP5972kw
JiRjQs5kSFx8gntYP3V2BuvIHM4fWdG7nAijoRDc6ri4x4JGQkzlMg8493MZHYa7
j0JJbdmmF/5tSD1lV2wizgNqLCQM/MW9He0/cItjca6FGHBhSx8bG0UaNvAxLqaX
EcVkfEFDsSsegINOEy3FG14137NI5C4YHLnD3iH5PAutlA1K6QW3cEBmbunJTDN6
7pqy6Fqqd9jZdwvlI3p+/rUPE7RD30vpmFIBJVPlSuxjaUYRfQ5Qz9D1RAEI3WRO
7volKjDF8+G+T2E1xVRQVBmPneJhdOy1Jo4MZQnMXun9JlkfrPlUxSkesrxYjf/R
0ZFzaoN9OECZGhscMINyX9Hcbot6sX/u3+RgQVzeyc5EH7RytZDvBrz6+cvu0Z4Q
aVmLNIdNgegFujhsLyXN3ii1n64m2pgqGQa8GzpeB4qoDL8K8jlBfXckp6prznMl
fg5E7RfCl267KUuAOJKhYJHqWXRi378nSLBOD8U+2CO9PX9VCQLh1WcOXOvq/qpM
bc5Emv3JzTWr3lqjyiftvrPgv7c2yS6gnSnEXWZPQZJdb0TJAkUegsZUTnm12ua9
/fAq4yJwEEbwD0/O6rDVhN4Tde/oStDFDP4KaNF8nfS8wSz9O6zcTRThhyk/+kMs
5zFyvwTugfQqWDciHCKbzS8z3vlQ4OmocsX1r6K/4CCkVhxG7+HaMYQ4yGvpJCac
d8+I6DtavVHuad1dJDYymfDq41HsPv2R6rPuQoVYu+o+i8X/E8laiTVE3YEmtaI5
0KjO3cKWtuv0d6rIAwX+dIfydhtXUdBss+8ib4rAnNQlAhbqnfdEbkU2X/PQvmKG
iZ1/T1Ikzga3Vj6Qw14bXSZ6fCJF5ZQ1QbZQUGE9r70FkcqBTiWvzWpczece5FBk
RaJDt8ALEHji/RG4zOb/xLeqDhKefLhfnendlcAHGeA82hEI/P91Gml+x6mrR7Sm
9a++Jf0a5SdriExYMsjri9DdbmDRsvC2PRoZL6viDwelzGS8NgUQ7jm95+BRz7u7
Bs16kApI1sWKzL7RJPmZsJIs/yGBxi0NPb42xztSUxdU/MgPmackU+buRDrGAODi
ZEkHJNIz+RkK7o85egZiwARNE1Xs1CtT7Z2+fFTvfvY1RqG+fm6OI2ZN+DSL/moW
18AH46dm3kqunNVXEWt5amswLpmcybyI5HFCIC1KMNkHeg+HayeIXFoIVhoyQ4E5
n5+zybcUrlT63J1H2/OIG/3a/6EvrmzuFi0efJi6or0+3N1M9Z+dwvCVXMCttIqq
kptH80+aiqqWEVgZJuliS5a3S3r6gD9Ra2kJRKEa6j0Xg7pRqtaIuOXeVUXDRmE7
+iG/7wA189ue8cS0MuYt6WxZiwn415nxDqtCO8dr6ui/DA/v2pTOPfhpiru1hVtO
FByEbTyutWjir9ZtNgVtqDkSfHzzLsC4RGgUQLfZRLBqh8MgHcCgFKxj35GdtLmh
EKJbxy9gbiZF3zxWmeAGNLM+feScPu+R33DdKGKVgeBjONMi8eYzQdAKMTEQtRvv
lRfb47k+MyDMzNw5BUsNREGKvy9itWoAY3BMhpCR3mFGN5UUeMe6o0QoWq1cqqz1
pMCpCanJgq16CG9bMGr0vFHIr71XYi90q0Q3VxQXgyRi+MFQVG3LKWkGvDUfTLeV
Qmb8da9zM8KRr0+u5wg3g6QfRp0rJ2gbhh0ZmM2dtkHNbRVx22puJqm7szDwsQa7
ihzyrAqdqZz1GRSWwlp1lUNZ74DJBP5WQwcwViKTg8lb62ZdrajGEIE0yOUX2zRA
uYvRvA+GPpwMMA+vOilWWyqP4hZD5o7DZEHWqkf/7kSthDHWjm6jSHRXmq9Bj67M
s8vllK48/xp6EmI99fvG0cbWvwjI+W7ko5IsO6LhOICzuf6HCCILRoQ55TXtHtKe
vgpziILBsWIASjeJVkFkGs4aBTn946rHJiSKPvutcyYf/xsSPcxkLGyn5/gNvn2U
uWZuKhD1zmczuw2cgWedwsb6JywJ9OTcXBhcm349lSfo4JgsSWoTpZzAs8dsYF0P
IuJ+Y56TEWYkJg91PATbfugzQ/Dczs4Gj4Jl3P77R0o2KRHamwmtFF5NbjD37Kcr
O+gjt0a9JYTRdkOesROyN4mzGjiv02Ib+ll+wNiwncmU2s6YC7gN+f0uxwA6gauo
70xA950rWAam7QUb4hZCc+7b5o/CfLb+SV1owxdBSiavi84jyLm8eCz2Ucja7OXl
4OHk+6OaVG5iNmG4/oozc4HwPITHo9Dnj++c16XilK8a6nzNvFObmTV7W6w+KVHE
FxIo69j8+3RakLKelsbDTyie1IfgbWKS0K0Lx6cnjUl+XD7mQwuZ91ee1Sxp2dnQ
uAO9xG+52OJwhYAths9NacC4Q3GvdKcoOq7QatTDQDJNKa4gBoMfm/7sqi8QLaUY
LBE2U80u13K5hX6qRLKtT+uK8gr9lVPQ/nXCAWW/yJZcFQcURjwd8cRD/DPw0MGA
MZlTHmsTml98gbIala5d5v2OULkL0HMPcTfy1Fbd3de5g942jXsXFlV4LbFy2x5R
jQMSs9miN3/272aArdVCrAaiLAO1CcEtPm5b47ARZMGOPgCUP7Mc8PzvUFFsx3yV
cZQIPDUtll55TCyJR2Pc0HnidcoW/j1kQuc84x4fKcYsAnj7HGpv7W6Qtyf9epFa
oi8zJVGqmCXMzcoObpVfjvpJcgXjIyIW6Xsn+sl0jWVWtZG9FqEGwr3Foc6UnaBr
xz6c54C1dCTRkAAZ758jAikaAAYIZMHlV8JsA5vdar2kBfBlxIf61weXYotzg0+4
mnnx6IJKi+KMifBVl7TqCs4wN1vNRqh5pRQo1HzlANUEuSWSt3CblVW+bhoY1f0P
+Pnnetp77JVPaAdLeIv31VtCczlRki+wVWKv5dESieRHSaN2Uhn3KCC8R9IeUExs
x0l5HX1KEQFY4wHMJwNgPDzrUu5lFJ/Dwe7Enlb9KSlS/Y5+ekkaN6rTyotCVh3l
usS8fsZChhJ4Jh20/SBHQPEr1zg8zUnRD0uji9L9pBXNq4iIQLmVLmZhgsU1x9Xe
tEX5uEZFmq7CA6vN7ahJi8r3ztq1Bz+zF7a2KGiG/ViKTNtSrZVMxlN4IQsg1PjW
vywullNyni2jEoKbcySGEZQ8iG8jDIzd/MdpTwh3i9ZXVfSUi79uVTPXP39EQv9I
x6EN7UmsmhwJpGEUu1vFO9HbtFxSulEMeLHZn9wZqb2Tz2uq1RlyeTitm6/wkEwT
awSQcWBEozhwO8fGYEEhi2UXOqHy6hXXXJo7S1okVfA0MSKHOlNToVvYbgWDsNOJ
Tfs0ctYcRtiwVlJTNAvsYtRadNcUfA1qEsKO65VLMWydOFvhJam4LQEW2oCCdlY+
3yOJRPQvS9PMWoVvNz+lqTObq75VyV8drBTztaOFTTs6zZygpITS4fJ8R2uRBMM3
w235HKSswm8zaLMKKh7VR/YXbWRRFFkNrbqSjmr663PwtjhL+cLShGOM8w9wWQaf
BhPlj/JRJXBg9Y2tmVoFcFF0pk63J2Jh69qqD9mihCX5rZT2nKUPGamKzqhliNts
u12tOGtyhvtk1gS6NUQU9qMixBaErWVcG7w6lCE6z8i+rNtinguxMys9sv6OvYH8
ZWZ7MtwD2/B7/DGPxAB8o66nJFQXE8Knzf2iSYQ0Q7zx8tnQtuy+vKDs5/qQ83Zd
cCUo/hkZM4NJEq2lJZaxhGYHEJr/dN9eFkAe1iW/dBkVtqgrGHHt/nP08+dIqfkV
GmOFrmlrsFnCyus6T0JSxRyFfibd9j09JlC3Ri4WpqBJAB+GWQunxgMlMklrZi5j
gRbrtbBRkEr1cajtJnwyNInKVgAPWf+x27cy71jSjA8VmcnON3vI2HjQcuAZlG3W
OjGq7HdydNM7FYQVEs6g8Nf/+g4sApBAYeh+JhzKZQ1KP8T72E6Uw8L2e5YGesdA
cJjpVI9zpKxCG7grXRWySA9ggGEMseHUClgYr6GjkakFuJXt76vaa03VOGsflPK7
g2VY/P7mqoVJXrQaOJuwAMa07Fe07FsiCsZYjZvf3O4CNeAM8kgalptUw2e5QpZN
s1brlPDRBgbuDx9SGC/bWuvX9dgZCXDwVPQclf+eK9dK4xWlJzAm51lXIcTOT5ZN
CE0NXXEZ+zPRAQ88/J8ligYt0FYIe+/fK5i2kMWL6XZoB8+j9vLUEIMi8qyGUbrK
CNI1TU1CpSoi6qXMRl9z/GBDo0I0u8lusTbxstIAlGh8tS9EyPUGsSenSgcgN9bj
UMJj+8Ko6LY7WFpxoMggQl8GCye7A7/m2rYKuKuoX9+3FIVZCaAEexyiF0X1kNzd
5D2HgBztnfYVLMX1ZS4mFtBdZWRqjn/ryHFVzpIvbvLOapp6p4j+H8xrkYODhKee
r9MXpNUF3VjjDA+0dFc2i9iRzvVb1Q9FoM+syYe/o7bQRSyqpiLewgupl8hcWoH+
0QiUbhajNj6MWATYcSwKqNK5HUmmbV0j4fyK4Ilt33p3mdtaPEY/YgToA/hi6Qz2
ZsdsKy5D0ZCD+B0eCmN5i69dYpA8/SS3Fh9vId3sMV/3dbtBOOa451FujWk+xVeG
GyTh2TMdl2fF8izsXdE5ObHeWfq2PRRP8rn8catoN1Dn9XTzu3XJwNrBAeld6gro
ui90oDdChzjtvD+x8CTSoPocwkwC5PftwpiZI5B/rL2iGnRupe+1jA3PUpEcGBHw
JzNWMEu6SJq9edlTR/BE8mDj2hc4UFxtX8X+QcjnGZ11NrvNwu4/oBWKeAfr9j6s
4R0o4vYPrRU74GOUYelS480wsi8cgoXTl+U4M+GUjgkrqFsWnEEP8rPQ7/lb9G0w
crlV+0B6VkAUzauVFYuvYait5yOGpCQmfb1r44r6BeDKq1msO6DoT1gYzwiG8vxS
LAb+pTjgi1K9KWbX6X7C3QiXukVRpw314JMYyL93QZd5WouO26LkFpxfIWePrDzC
p5pVjWgX+mHKRkS1wbdRsH3WpOXESftw9WOcoBwLtGqx1uGRia7DtV9PIzRwiHGD
5DBqpby0LLXbf8yoViDIDmgf94n4d5b77ZMUXjvCdrGaPnk0zOHS2upVnQC6dhIP
ZbMsv5DyvlKfzJJ4OQ4QEX89nWdKt4TqW7Cudh0DseoD+syY2R/uSINosQAQyE2I
YGOlmN81QEaozAGIxPM9i5uQE2S2lwee6XWU4+aMFeTeSuYR5kQwjp8PhMGvEyKQ
sHg82W4jYiYkodG07bBvlp8K5Z7+QR86usUyW83+Y2ynTM8PszXgNP2BVHwn6qhC
Nj4hr0+iKTQnVlSdWC9JSs0B4DDNHXjit9C85lBLCkoox/so85yChFP2uwjYSn0N
gmHZPe6EgnLoQisLkrnPdafYCgWtonBK3eWdxWwlLFZ4pzegxqiGGFSq4xSSsBLF
aRJvblAIr8HA4qNCfvA5bfkduzCLztQLQ/fN2KiT4DEfSCNtLfi6Y8w4AFBkQIbJ
Y5VliQAhYfeDyjsBKF2+4LLkAR4QrOzvWa37mR1tuB8l0C5RdpS+xWV4wkq9HL3I
dsYserQ+sbK+5Nfnr90z1MIV86n0zmmsJLOfY4rMNA/cld/I+43QP42n0Hzoy18j
KLy0zvA6TRW2Zx5BMnsxTKzYbESNqjw2AmEh9cGFe7B5X6FG0OuGpoFxC65rumW3
MAzoYxejS/Ah9lcz7egSC4LDJtmIUyQQNUs512w4YBRO1zgWBl0Wuf7e0Jx8sFa3
VMhZ0RO1ZHzG/0MoDxqkxG5cuKCI4k5nEkla7Tx03zVZgpZAJMDM+DAWYkYZ3qum
wQy2F5s37PmDDtuTdmJeS5OpWbAMUDnnGChZQBnBRqZE8Q4D7BIPWkrJ+Mk0AZR9
qbXwwdADBeKZTzalmYHxoFhgvsrhGnVf0Sk2wcf+AI42/aybyqrYBYl0tY3/D/1j
hQ7snERphB1vqnWSJ/kNSvEn4Dvoti3u5Gn4JqreVjDbNcunSfTT6B2gqA0j1fzu
vYLF2TJM1Co5oQrYCQnc6r4F3MfaLQIgMjBU5ml3yv+9zn+qsia6SAbi08gz45ar
uy7rTdyGLgepOYls4O5uGIyut1Z554rb7MGoRfzFYNTSst8eZ03mW55ZHKgRf3we
req/XkY/r8AxugpGvhC7cg4lvQebg1M1nrfvy3Qa9iFmnxIqQT8I5WUAGNnKS1q3
ZilcDJFzymEXqgcpuAUeTKtRro6Ztqenv4GpfEQCbXFuewPuKuVWxeChgZxbsmcj
PMtdx6ij9pal0KXHwDJrMu+S9v/QBTlzilS3v8udJ00Ey11ndmA4A4SD9fUk2zC/
GXzARTfkrtSbM0CLa9qmYzK4vrO0Nje0QjypgtZ1fe9yVPlND1+5J2IWTXyaVp49
YV+ZE7whwrG5Wj5j+qI+E0jyYz5QCsCzFh0lhpfNGabYvkVuPia57KQXKMZmTD0h
xKhB4DkgXjmMUs2tQdvW8pvAERwNkTJ5ZFS3NzoBsfEtA6ELiF5DO8ue0U6xFvmR
i/AZO5agiiBBf/DJ45vOAFchOn1nUgMnY0ASgBUdMxMGLnR9ZO0e7lSqtLnM4lD2
RYd6YLH9jL+/rlR2Kjz6swEv4oS+OcSvx4t+BOoOY+LcTggEYL90DoYWw8zEUb/3
t2i+RXr5hopSkmJp5VqWigf2dIHYCfWacIYuKB7M3Z76xShw6fS1B9HaYZUeHB1w
d5JpV9YJQuMbLnztaljCzvc9mz6fPQFuBCflGH5sd6u87mtwxnYzEynhJ7Xx0Z4m
3dsu1jiuB0ARv+DsL0fU5erWq1afuG6sZHRD0BNc34PorPSkzYRBXbIrFo18PSxv
dkgt5Vlcofv7vikhKzNOe1YMjFWfBHutCvufiOakVbE0UUcBSK6NqxvyNWaIFr+6
B6MapHjZMKQtC5TpwPgdWpZDzSKlumQyKr0kbBDYnpV4cLRmTKVvL+smcZQ8paMc
BdG4uOI5jF8RsmJGWmSMpjpVl6RGmeIx8DN8R6ouFkdeCODloCqyGOghm3ir3q6r
iPNzQB8eS7hnmLW9ytthONxFsY+3Es9CsgQ0hYDkj9z6KdgF12bswHxwJHRVOg7H
7PM8CGE9bm0BfmBDXQJ/LPGW1xyWx6UGBPlOcN2cvrNw16ft/62t/ZrmQN0Y6jpS
wRjo1PqOdN9IVcKhcYYa8C3wdV5lyyc7e64jF7Vs0Wn167tuOVGsPE1r/nsWEd5z
bBNQuMLftUdJMe0wgE4uPclrFn0FGL4f7sfCt4nmJ8yHDsfTFxiAP5sdlWltH3Ms
WqLncJ/7AXqpUg38niB77WT7mV7Dl3R0Zz8LanXOdvkS7O5F632QSlnamnaej2bk
H9peEzF9wAIYlChIg0Kl/IjVf6JG47STAzbKPo1Zz9JUslEx+MpTlE78ZuDh3RkG
a0BHR0EbnM28J7rm9l7yoO7qxOZgINbxSGSrhnU4J8Mpa+7kQ+6EkBx6wlNGDr4Q
YlQ8pFhTfwLMfjxj9SplY/Xj+witixGY8B0Nrdb9gfw/Oxt0VGE04avxNdLooa90
Yru5we8mJIdtS2h7YtcJi6rCCKy0HiWC0YLs43pMkzpXw6end8Be68GMhkFu+oGl
WRbiMKG3gUz2ObcReYQTviWUoBWmKmFikhbRL3gRmNBCIZkYg2jXsh4SxFMLaOeo
NBejzsDyL704GpQEVw3ciKFqACezEEimwr5Wuyg3MlBNDVoQ1js8vqiJ33JQml7W
haIRZGkgNgSrVFqYnNRxSHooJM3XIHjvFcHXsp/nErS/iTH601v9KBskq+shpy44
e0EAeXZNLGKj2k0+JcTPvwZkMKiHk8wjQG6BZIt9QAZTKA7TIoaK9O3Rj3ottgWC
QNr/RRLk7EPguTfW20H9hPqu27yeCQ0aZ1ck0nQ1uAg4zV816xMNkPYtji+HWGXg
ijgkjr7dS6P0/uUKTd6QzkyxCsiTTmKjGc2kKBjUi+9UmsPychGFe7jDAUpTe/q6
m9lCwgo7WU1CAbCGaYzPrnPO87frCka/iFC13fhWpzj6IhCJuJcfqrbaI5vrkdfI
HrTlYRHuTEECO6DHy3XNKL4oTLFKkx7I/zKgf9T1teiUhwdKnsp1AsRoyF6hJlou
pCaHOKCY7+R9n45BZnPNaRV2EyM5zSKbSJVEBIPMaLWhbQRKFWYLBZ5k91vugFcl
1kkYrIvI4dFjKFMnIjX+yVzf3JMKJXvowgfBrlSh6y2UIj1gn4UUYm2D9MF2quOv
IUkNNMctsfKeEKvL7CdCZwWxAySf0rDoZ461JL+UEkzwQyhsKQY6ruH3D13+2C4r
VD1non0OrBmcTbyZ0mQDa6YHwX7Vv9euxEocuvVa22zrj8hsQX+7au2gJqqwwsW/
O4XbtwZJ7fVKqgI15qGP/kgQruuxonDQl1eR9BhMqmLuSqYa1wgq4t5GPFsEnT/p
6SjriPg3V7dB7akVkivzCiH6MUyC5us7puRRLl7PBORIeIk7sHoJoxZt8My6M/xe
gSTLsahwhMZ89tT7dX299UCd5+li04OOwHmc6MYXqsNWHFNjbCJ9l8XNEfVzdX7x
bUmqsLQqDpf138m3Hm/xcytcVDSQVYvn0hjcR7HpV1Sn5+M0r6QLiceZ1h5LKY0x
HoPIWMbGvG4evkDX8QiNN4XNxawiJCyYPkydtgV2zJIl4oI8aTgHOOzmCvNsFdJQ
+Iqe/Ag302WzNtIlcoBYqnYIPkwpXiwCMDZKAotU5AuSgdBPmTyytkHk4Nn/7uTW
FU5OcftTkAzBnVqFCiTzvGguxVw07UZWsl406qQu3cCBiX1CYxfLKMCrrUyqevcx
E/6E6RnEpE/mq/e1JRQgyqXER22r1NU/bRg8Me4uoZsC++h4MdSPYmCeZZKA3fv4
qOW697yyJWXE04GxnY/rKxKONS10D2H6wo+hGnTzLq/gyJ+cNMu/vq0TLavWG0Vk
02Gk2QuBZ8Y+s4F/rO1mwX/p5dUiHgvhshCsZ/TF8USa0+UWkYdWCambzHHtjazS
mszEfynwy/7vPQSijKhiXfvgO937HswzS5otbZNkYnB9LkEwREgcIPLgRH96Y6nM
XiYDSkF+6jqVA3svI7Bj+1++yAA53/Jp43VKK4SZFUTHgmHMoXfxLBKhprmiN40t
DYZmoRm3ot08/Tv2ib9ekmq6MBB72gNs/Nd7loWCUPUZ7k+C5SlSIo7DdNjhWIWN
Se5wYwRXdt9zABjBqCqamfBfX3mZd1nW6eYvuEdwX10XUYWbKOVuDBEvR4NWJeEC
rORJY1+grP05qOAdpsuopVTtb8+aVcs7jrp6PWFpjITcizY9uKqz2sXKy3SRQyEi
6+/V7fAlQIhujweaMzI+677LuTgLuIl8W8H3s8jTr0kMnvlCTcuMhhHkyvzZ/hQn
D67BMAfQ7NcZjBEdQ1JmJXbjwlp098YZTUGdHKAlPBGG+/1Y90RymeRQ4JUI0sKq
+jXrnQCQg7ob/GZYt/FlgROwBKsRP8lxPsp9K+KtAyoUujqSifjPhPJTsYKMvvFM
S/TuIhVsWq123CE6uMcaSqBuHIOxxPMyYQUgxkYAjkN+axuD3sh2rZVyo8ifvO9Z
69b1jsgnYENEEp/K/a7N6LZqinWaA0HKEG1I9vVmwuAaWiw/8wJr/nnXjAAqvJLF
SqYoV8nOELgOn+1fmH7YxrRvIwsBmD6ZCalg2UjoOYZ0mxy64+ciIa6CACDFAH6d
xi88uvfOYm35m8u5VEsThtDBMQyx9LYYL5ss3v7BCD/xjypHKD7ULuhh3BbadZLe
ip/XnRtI2VhsaYNctxzmbRF107sGgPCxo8ZhyBV3fvCQ+lzaM01kmQjKehIZ9VfZ
WZsrnn69DSnxPl18cz5GF3CeKsKEKBdtBFYrzx5K8fsTqRcq9lg0opjMnoG45wnm
P2fs2MBKdAvZeQ+0sBZB0JFJgbLoQnLdv7WeKOd1qROBPbagKPCiuG8J/CWNemIh
l3oOL7tdkWWA15TnwOV4CfV7oowgFwsCAJgmMRDsk6ticiu/PA43ILpgfQZ9NjZ2
E4bqRLdiEKMzsylaL7xUrJlFEysCRtWDWQ9w4ByhiDT4+R4XBO3RrayFT4xPfUiZ
Na5gCqSU4rmpwk0SdpQm7mUZatMHv1VZfzRG4afwPDa25S7aERivN8UJXaFoa/TN
Fl/LwFRO3+HUmX+yoFyo74aINz35vqa+93oNTXz/RNGMLZVu9WOdoEQOeVDqhJOS
HG2dbh4QO2lss6D+OTYrhg/58+1HHndgQNxmneApegC+daaCPD4kCrSRKtalpVSk
AltyB0gvdJIiI0h8o2HrUSR8AtSO53sVbC/LEy7Az1/FxJNDGdw1nLKyvZsGiJ1W
poLukBmA3xrEj9HUT1r/ulQRS6t+zj7dObovXh+I2YEEaO+RjQG8mn4xb6bp93m9
bgu6kAIDdR8J+wI6d+ylrsIHZKrL8MpHX3FupzC7J5DGnhq6TaUxq0z6XkWZBHzH
s6HkG2KzswaLc6ZuzZu+AmvlHY2k5Uf9gAp0yEOUJddX9kt/7oTsFtBicqBwvW7r
kfELZX/Kq3yj7C1aFxbIlUioyzkeDdNS8SGXMkhRBkDszKSU8XhuK/TRmqiLvrFV
N4Bg/fZLCPWKIoenkM9Mu/D3OBX73L8VaKH8ZnI0lGkBI8s4dyc+oDdSGVKAYPNz
WXi3/qloJyyhV58M4mnDRx95mppqMNUZlnPh29yozROqGtzbQacUCtNGLvxBkYG9
nuyxS/17TMlgox3rnoYfMf8zZIprb63Rj4IGommr8QsCccS4G10tcT07YwC/0s2b
VTJl7FZmka7a1Z/P1sr1zvf1fxoEuQnbPNIRbWMklaDA/qGV7OjBkYin0QAMLPwL
5SrVWzza6Jaf9Zf7umI1BmDA/Ixac2wXVDhsg0IXCY1/Ce5tRlhuwWDoChYYbjTJ
+PTJMmrUCf5oHA6DkYyxv4P5bsLBdNmLZy/x+Lu0o2poXlQGDOdf7lVneH+mV4cU
blu4IqDbmZkjSuX9IFHInDKdwD7WO+y8fBZemjZ0drsIrDT1+kPahOZLlzsoiYgI
lY539ewClVSf4ZxIFWE7AMswsEv6YGdbM7cA5LdMwRrDQl+oLGItImgJzD7g4UWG
y8gFE5q3pW8pLWyyIwHZT3w8z5qC325cFeL9HPsoi5Qmwj7XlWUXX36R7/GtiKwC
tMlGhckreCPATJL9Ma3WtKYzP5e7tl0kJ9rsmej1GTb58TeWPsqShLby8uUg35aL
h1uDIdXMu0e0AvAt7yzsWmzMVCTx5TDd6fxs7r5emeSls1vsxcHvRtASjHx0K7Ky
21fAybqQCrcN3wqkZniVGaOryTZ8BpB2nTADrc/0L6i8ejbeBwjLhxOtnWYIld2K
tQMBBMTeFrLenBpnKKETnNq9+qoh0QPDyC1s878bLs68i360gCyLF4ggWjZpJ2sw
ilbJ51K9WtWgUttF5TLllLAOuZ3fh5UFM/45ZjJTD7MiHorEPN6BKbDM9KfNjgXq
4lmVYd+I6fGUo8IGCv7WOwnYBhTtpq+Cv72zkb8y8JqIo2iNEufIf6OLp6Ne8lst
z9QfKnTNG7hW+c68qYNs4+ECnNwOAn3vmHwhMW7E6FozuhIEr9ILZ0l6a2kLkFRw
yg0T12PnVszAwYXFpGr+Ni87NFQAa9sG1Ns2e+7AZ/0VB0aQ3o0ZoBFnN6Y8mFHT
cxDBZbUNcrXJpm3XA9mDvOaB+hQHoXyuIFQBu4FdxnGVS9ndu+vCsDwVSETteZGA
G9lS9FSgcNvcn+2tUH0yqrQJxdVq9Mkjge8OgC4auAb+h3UXAgTIa9OLJSEqk2F3
RSubRhG9mAUNH6iceEVM1K3R5LXN1tRDw3G20K2em90mMKCmxzFWeYVoqcCcI1rW
cAZo2ToLosK8i9JHwDtvEL0H6hB/DL8Z6j8XRHsng2u6HN4NWvDCRQ0nK412O2CK
7elVeVvx3yCqxSGMwmupXfcTlmAAQeCupmiHYSSHv2ADhtVdoPGYstd355wnP8GN
JtRYnRbxw2kDl9r+gZGzLcdhF3G/hHlhmxdI5AiKBtoeS4K8Bls1ss6GpUOSllGw
VV44hT+Rz8CfQCZUU14/qA6lKfJV4GKNr9MTQ0ih/aI3N2pmSIlgTQwsxWpdhhEX
myGNuJ5/QAwErUJJ8uEu9Qj6PPf/vhVOYiJ7iCsICyEgDRo9I3XraFwYk985f2SS
xz2Tq0imYJmM2/Mszy41aAcL5PgF+37ZC0zyA1JJFSm97RIEg9vyh/dJ2mtV655N
7sLDidK7ashGTGgrO3D6V2PNShnA43VuZvW5htCaWz8eCGz3cBmYpdYcZ2EZDNft
xp7oHaP18IDKTqtB435+ylvAFc4oW0c8lc1Q1LSXsP8HvTc4WCm/Lnplm74Uf2o1
GN6IiIHed95iXtRi3fI+GQj3XXawv/7uEj+yoWIljs04Nqgy+xr5jonYPw4fGFiK
MSQTkcDrvssOe7A7cvL4sz2+xvlYW1OPpx7jfuk1llNcd/moweRvOZZL+Vi9wrna
rzddito7OAJIIQl5HhfcXuxzlDLvWmWDiWNYHzHTCjpB7TXyYb3XyYDl01JN4ZjM
8aiRwja9G3VXwAufN2nIurVLGgYI86xlTns0R1g5KaVf0qivMs9VKhTYXwYuG7Q6
lHwdrEcAviv5ITbmhkxI4e++fYAf0zhJFModrCwdNhm5UeCd/3Ii9VE8pu4E7qfB
iIFMo6QgInBpJdhkSuqvOJmHT8W/D+ZYAnmI0qcj/HszUycasB1uAGdDvvrwe4en
wUPapmfosqvuSMweLDHv0XY7DzqZ/DiTZbRkrc7wfn91vyrHQTr4fy+iCaNREOf3
epUHoZEJ4KrkDqSht/OLQaZnHOy49WcR7bY6lEZ8ywT4KuYRTBsXy7x/lom8kRDI
hY6jGVIqj4yvDAsd2lxM0ovP/p/vcPE0bl7r/35l8N2ZoFwWmgc+c34AaWYvWdCU
UUJkMblZhMFr17EzIaeY4Gs+E6ZKB60ppk002fO0eQVbn3jIU1xtFfGQ2Nv4gwbS
aAOO2/zMX+1FOM/SRJjAsYuozThjh28YJEzb1eLuwrV6lFi03I01O1C3fuwTHWmB
7q9d5IRbEM7u183HRm58p6ATc+6K20RJRCCgrFMh5cTuhGq4OUXvIi4Ot5uQp9P5
P3BiYsFZDMT8EVvNSomeqriWTqo4Wuis1cg+74SojnVRY4VX1/n+KSMTwzQRwrnu
pfKOPVAdRmPvIQ06pbHLmgYX8jvCWkabpWg90q8MVG89o4lRWJSKCxcbu/tc2mIY
BYLmxnmDvHHJzMt8IvpP9nb0YyetFj2pIPbuSdbVOhXsKzJItQuRnwijwvcHPx5F
nISbhYEMfwhXnTQH1CDFiYGY9x/U7PJ8nKomt/XdRmoXYHC/IuqIeFWyxPSbg08q
WuPN+oAsLM81+murM1vQjtyO0vSpSYS70f13SyQSzUB1ICS4FFjDRT3NkR4uWeF6
JZAJ8jbbpyKQY0xX096m4yfx1d2VDI/RutpozRsdTJ0a6Bt/ckBl5syxvZ9+qyjY
yAp4hz/Lt7Mkj6wazwS2apCYfO5OFhf/+7khpSBr32cPW50dpEGxc3QSYMOy7a8o
mJIaxisHOGfXlVIYQc6ryk42gLvyM7/YtrcHXN5sALa7lcvQMkq0+evCWoHKPNto
0PQQ6D/zF9mWe1JWC17APXKkwTUmjtf5m4a1jmFV6OH1ikQINYcQg/KyX2TWcg7f
fZ2/9+rGEqMA4ogCMyMHyGJpppEOOPOkt4oAVGzLeEblcvdfgVeDPLdslgl6B07i
1waRiSDLS3D7AhtkzqMJx++QwxgeLJgKZH0y+bBFtKum6q9UbOtZ9DmVtPGVsRfT
jA5mioslK+N0n5vQD5RzzsO/09oJWe/49tdBk/p1qqIbth+YK5uOVMD/0zsFBlnl
ZJhFIMhcuKhWucrPxIdIZzT/z+s/PPkS3u7DVmHpy+DgEwKYP2QJaRAb6kJl4RzJ
1QOqP4/pb+jXCXWNCfZPGVQlpT5kRRn6OeTGcXU/U7fWdfeAWVCaM6+5t9P1Ysei
keF2oAhAO8aeoAJZ9XxrkUPrXjkgf7OZrLSv4wqbcnceCiSUsuz71OWan1JMXtdV
2OPbqbyeVSb4q+FQ721mc4W9bQaMSPBq7SoIPq19mioHNN0FRc9TMv2UMU7Ar8cz
XMdd3bNuSElkLrBrqhEu2qebvP6Y9PcFBlOM20kuQnjFDRNn/eqjbCUH4y3I0pbI
uOFclgohQveGqdGtYUCf5Ub+CfKvSAmnOM95O21MBwOcZgCrqsbN0SLJ8m3QiHGQ
65gl+XXG3rnP+bIl291hVz91XNwKrGhFqTp5abbNHYw5TCPxNQrLdf+G5uC2XFrQ
aLm7RFe+Sa6pmRM7gGync5sghdEgcEtA75WmEE1NC7N/MKVx4qWvqvCahNHAso9W
zmxZQQATcrr0DuwHjioso//N5jLYvTm9rIr36oEIRPCkCdBQ06ZPOcfYMbuEkbGd
mFPklLrNjZYPg8/LHS5ewiNffHiYY5wlzxQ9nrU6TpDg5lqDBWyq+kj5U0aQlW3q
QGq9v+IqQ2yxR16AUFM84wD9oDPc8bSchgEh4FpzLMU+6ES8DVhsPBIbt0wdLk1e
wSkiImklt+cU2XeN8yrP3zSFUvtCn+QRVxv/MgmreroZwem9Q2WSHU4WUqglScYf
oWWRp+8NMbCpqEv+HVxjGjY6tb8h6p8us/Nb3279oq4rzmrWogH4F4DsPdFsDWYk
03eOjKRhZzFX3Nf7Jkrkj4idUFg0ScMBCsAt0T6Ssez9scvAeNN4pS+PnCyV30dG
67M747CHmfExnAanpXAKZyYAY5D7MHK3jgfCcG5TPB7v7Ac3y1FHkD/jnA4D6XyH
1bVLhHNYAW9AiAdJ2B2zRp/rLVxUfuRsmqw1Xit4XOPZA4/fHro/XjAnh9D+uHhd
BoxxlTHcWDvna7NFEfidcnXjMK1Yi6DQ7JO+l5giZ3ax9INdlblwGx8WMsdC2e8x
9MsZq6/YXKHEUw3udXTZxL8m+CTuToVQqIH0w3PYmPu1Xkf22R4ABr1c4HZYy+WN
on9BQczpG5DsXOXyOldglRo7cizvTFWHcQQExwUksAW1Lg2mqGDVDWOOPYaoNTYH
dOtDBL58HoUX6kZSjK/JOPYobpUxtSUoZqyWxwNch53khErfofkUgasT+dBWQZNa
4BQ/Q2Y3+uBNeONdmzJn0vK0z2MZg9NgbIp+Lpsl2iROquq5ZxSGVCU/IU5eBCXO
+rN8aWZSW4RfbBoOkcWtuJf350+mUbSOkTfnmNJldGBMNVwH+1FlelYzGT6pqfBI
E8uFko7rjZNoSMSohCWxRVhdrheg6Q4bpJVfZAv0fy57NSviGFX4JA0uggM/SmQ8
ztlXbB3DGJ0CDr6a6Gn+Rzs6C5haC9LCLe9ZfJlHzpXEVZbb/xJJCjVvxjBXfhlC
uxm5HZ+frtGRCr2JF0vz+lJy+v85mhxZvmCIz4wHGo9+hJOqnIfKniW5XWhU+juI
8Ju4bKTH9Pn90GvrWvJp4a620ZwhjdJPykidiS2VjdqAOnpY77IICJGOQbs9IwUI
EfBgM4GmlFwtzgVIRxrIj1mfcL7R5uk+SZ+fqZxxgLuzuL2WXfbzi9nOkvUZo32g
nuwzd+N7H8fxe73Py6ncS0OgvWqcB5dKjf6NuQZ12jviEc8xUEzrOnVPm4DUyLsF
/8hoEE3Uq9hgGRSfNT57J4/+miNHrFYqPymV9L1/e1kg57JklU5RpZneJO9Z4++Q
3UxetJenpth9zv6evoMYvglghW5YD/4/2lPy2NUKQ+YnAdokXwrE3UTW81XNtDli
PDX1pg8J5eDInpvRYnss/tho5vsJcrInMPjABPIkctY5/82HieGaQOgp9DQGpMx/
CtAqbl2bzfPuVWFSPebfhkpx+8owSXFnL4CV4NtNTIWImpmKOuJQg/mBuOl1NqwT
WMKEuOPN55KFH71/5lHqDeSSyIfK2IIW1pbO6vQYbjqiafAlU0frDr+YIdp3jKH3
dxMjH0u0Do1d6JljUYHNTDvMCVqwl7fGLUnpbpkzhxMDR9M8R5pXmUaxMhiAt+Ac
cQtHG436wD7ldub53WVaMhDvvyRXlrhvyf1BYN439RLnxWWZeswlgphYkldW5+k5
jjlBGpX06XFSbcQmrY42l5hVMy3vKmCsp3L+emTs6qIJaRD0ikITFn8Dt8B8eCJa
6ZKsbPT35yLIFna4L7a9nwsKI3vqAQB6gbobSHbGGLdl0Hj6NfE0a6pAqtwHyXOy
S1FoFFVzOdSxs/uLijWyrfP0YNIwEIxpmMPAezcFOSvSbfv3XHpf4NQ5yHYzqkaF
Q+mhdspZyDtlLzFABgS6XUBfh1znIgSa3riJ9zrnFTTsqswie7rkowvzoW4kCaOW
1FaKhF4ZxFbJ1hlZbiTc969KazLMF20rmhjHzGawEw71DoVLcIUV6h+HfdMz+tBZ
YuN3K6gA/81UXpfAGJqCU9+yofgo7BE9boFmVeEr+U6U7oG5szHJVQQ1SitbbxxX
M6JGirIT4oZB8CEyUXGp0fHtATv2ab0J/WZRk7nJYLWQzm9gEOgSncfnc6RrCAC6
2IaO1Sd+qckEtYFa1QmyEdaNxQn0eJ4MAIPw7B/Xsj76Aseh7RFGflyx4B29Rqzs
/rDXlowsiV0lDXMCFn7d2I3IMdJs2SUqtsx0Jtx0W5xHge2CT5LCmk9PnScOnWY3
SXTvgfJYTxuoryOlmzJSMzKdMnqY+vf0QxhBxhtU+44MVTiJmxSdrXqECECxkaqh
Ws7r1DJQfCNe9CnSSTwpsXI5SI1LBt41RZDShzHLRtWufA+bzNKZW32paiSJNrJF
69BKywWXuZIlmM0z9kTfxyfFfM6rG1S2t49uw77SFJ1qmMzuElbHxUPr5CRxvoDP
8vSSrQUHqBMBctRp0mdlKF20mhOZJjnVWnHx5MDSVIKpGhit2I3qGNbxfu2VFbuC
7vQvCldGhuQAiTfYAxV4ETg574mmB93ox/8wuPA7PCClw9HZ79soAczW1uD7uWol
XGtPJ3UN8+FqvTbbrbB/P08etKhTcDDTDLl6ZxTbuGktL+O5lmEX3+dAIzGuvF+o
OjX/JwqzPbvEEy+DHQOSeIcceuqMEyHDGWOlYDS37sx9qHq1qkCf2EANZGHTJCf5
Ejr7z/p7Nav/83vCOUnrtG8TP5o5YeGpAH0dwycNy58AFZOmUkeY7sOKM1Sbf2Vw
62ikRQHpx76Y5ojVkOv/WtOFJkXl/iO2GACriWCUU9LLlU+/gZJmPOq2Hg0Q7mzw
CxlNtlodyVAnSIEKsxlVQufOxV84Bn8/EkmwuoZmou+z+eEJNk5sRu/AudWkW4dg
ijz7PvwzHYwGQ6Ee8o7mREv9ZBE1AKr8yPQSPpX7ALDJscCkGWecnaVNBvIgoJA3
7jGfUE6SiQK7Rt9a/RcbpCOrg9/OUFWvO3YVX9/lBBNkWSCN5E77vJp5yA7H4HFA
KeJ2Nxghew/o3WvoMnWtBHdXAAUmwiWJgPEJPMW3So44ERD6Kl79Df99M5/xwQWJ
oKyoAwzicmBHgc8fZAC5/zh36cjYtMWBvfPinPBLJYZdNkp6E+bC9sM/fHEzyp9J
ESodeIXTS7aaavwEaIQMc+K0mTjrHQWNF+f1vxeM2QY9+LewGPTzPCCbthkYCJ8w
7wfDKP7Vvs9Cw6I/rFUQGIVwHfvWQAwbVpP0LfSWTMdJTnuTxw7wdhf5fSVh6DvP
tZ01N0cs3B4XDpvsvgk2XKzgS+MQ5uxfgLkQ5W66nWC1F4uK+I1QtcFia8FICRJ2
YWG5pxWWEgYri/Et4dRFNZlS5VzM1Wo/khTs3i+AVURWUgRUQAuDR95XS7AlVXpE
mKVSCnBEEYG4twQIcweKNzWqqEsJvoNxCCcFVqe/CSsx1EWkpEUxt08pEzFfgrTV
/a1Il/d4SJMaue3FNOoxfqVaeeQhWQScEIR1twCLBuHCAoOkChgBPITjdrPQ9yhB
7ooBiOOke98uKRjH65qzDiDV0s6Wu5J3Ta/WT6sGRu5PW3OeiDLlA3NpdTvzvZ9H
r5feZlbFFhNQmdRddHXnMV6UDt9BbsPaTq8tbOtILdp+hvPhQQ8BeFQLxOtK1glx
CEzsvzXH6rgzx8VjP7Q/nzQU6SEHh/kckSCb6UNL5Z3MtNU3Tmw0TlP3xR5Y6zIG
w1gMg5yFj+tJW40rBhs8N+if4Osa8LlBpDpqHWkpr0Y/0ycyw5vdoTx/9OU2n6dz
SEjkrN54byE7FuMWBfbTlDU6k5ZKZy3mwWSaMJ4q9v9uflk64q6zzEcPWRnMPN3z
hz0OttQ6kvg2bqQQ01ev+ycOoJRw6SJ+emoTeYMp0plAi6kTbqTZGeBG0WfGslbh
v3Jx2oJdCtOriZ/TqYWsXeEECfTQhOsHf8B62sBz0dbGUaLdAglbvTze4vA59gCX
ZZtSFTknvVAKPzSQSWMnYSSE235AL61t9AxwIYneM23Yzk7vMUx0iaoe3+fDRq3I
DmjGu+PrRQmF3BKqgEsIsQg9dqsOuffGUuM+rwKpnqOVv8JvSEv3Zg4ucpJDm3yx
b+8rp+WzokJ1Fgk3IzFIwcrAqfwvfIFX0KzitxSUcEL0xjYL2gnwe2H88D34RNRa
FpD2NOBSfg7d2wZWN2oMv4Mdwupr54vWz+5Ayf8E+l0TWU9/fj+Ke2633IykEZe5
WyWoM7c7ZjLNUEF6kugJR3RuggPVDlZqYUNko5TyjiHN8XewPWubfWmIvhfMIRs6
cm0WTxVYBJuiD+um4aowhczHZxDDA4yamRdcTc7QEnACa90tgg7PcsvhrAnPk/pX
jGmyri5YGIkjUgDvGWWBpaUY8zbfcncPX0KVMflegxfBa5geIEN0qIuo18KI/3h1
cPW+YhKbtfiysZ96zhW6K/yWscaQ58iFFC0EOvV3o1KncfXFiR6ZIubiaccpBxSb
pqOxNtzcH2bs9++G43weRpnpLEt9pzgNZL+UlbEHeoUR4bqFrU1rR0FG1NAtxKBt
vUqveJvRpw5CwQo9RbC0tB+8dqT9FOX7QTQ7s7WgDJ6SIFRYke0lKbqSK7vuJxG5
ixlWAS9VQ57D1UfMhmpp5pn0tBEOb/nvckkCNe+cHvYD9eXfUZdaKR3xDbEUP9ye
P/OEYtAlWIbrn3Z5/kvg75naqnwtlO8D+qTgCIzM0oseAbJIOPskRoccGUMRpXvi
iMObeBLXUEJlsjYae6FFmSdoB2UccTLAYomMdsXSPGR30y/vIJ94EYeTkRHrDdws
n/piCwbmSEU5CrfFh5kyB2/rvpIP9Ce3nmFJwZgz1KRZ0qcszQYWhkOazA5Dee/w
xBMvaKM8XpEEISyo+yFCwWxv2V75el1pNSL0FEhGSOwWxE0V0EytbALPqLFIZPCJ
EAJaLlbZBQ8a8mEgBfGaY8a8HESXbiXMpXEMrzj4m4EzjoSwBaT343/fKmtf4OWg
N/sAd6OnUDYXrj6IJKCgrdFj/5Al5IrircgT2Dr4zHbToyidsu8nGwWxx0WO0VU4
j27seaAEaNcVI9AG3Z09iifYiuZ1Dposw46WR5U7re8VHu7X4zJBFlrJxvN3uw6s
TYgnEARVCGvu1ttFAj1BevTwokzZDFImIlnkDTcdLxC8PUpd0kejwN/Z4P0grBSS
CxHDXbbCCD34GMlTGNo3EOYf6Ex7S0Csxgmmevu9iIJOlmdlBD9Y/y+AsXM3TSyc
DDgjhaqYY0Hch7+b1+FaEOY5sFXZ3xLZ4qy3rwLXqOuCfBmVJmNO38gfaZkZl/xn
svz7lMxcehEJXjhguZ4oqxur9Vz4A66A1p6QLyi+HiS+9tIjWdgu9vSZI3ey/U8k
6caHLTEuD8yJz03GC6N768UHAjU2LnTpG0776dBEQCY5CeXYQuuP7bhWoKbt94hM
ZKfvHkZox/AyYVEvHo3wFjYqtZwB04qjmSTNSJwNPvjIiGs7fiG8UzS+8ixqyFTh
Ji8RwQev1zbhPxw1ECrrZkQPGLmtHrroxJO01qOuNPnqLgUvyO8KcSD0VtmSjOSr
VAw3GO2OII60fvEPjYTY4RdVINzCnFK+Av9rh28vor+qy/nvx2BiQSJE8QWAuK0G
BHaxoro31u9IQzolmOLey43U4C3d5P5pcecL3oAKmtW201V0oYardcZDFR7B3PEl
SYX7lUd5UI+o1iePAt50k23OLFL0JnfuIbkGEn/m1mlpVbKEf8oXa5a7nB8aXLA0
fA5BD44HFx4BfspviUMhU9X8GJrWogwy77ExVs1fS++xJZCN4jfiIeHA23h6FcUO
RmcK6M5Qrje8W4PrsBiJOXkfp6gjVH8bsZyyHovoZmpJSvSxjyWCfBC2MNtKhy2T
o0juQiKLQqzUqhWUKhoP3tkZKphrKM/dmUqNTvVEMBC9JGP+mXcIpO9MCkNMH82s
uToawVH+zC7SFODuQ4G/TmJjx/Ahd9jOuyizLAxhFJ3zjqH1+Vs0UzrqBPIAocyQ
KQnPlFcIHE/e3gEsirfLiVSa1Kh/eVANKN8djwjHC7UmZ3sPP9PPXspMGPTHng4W
R3N+Zz2rIZq2is8lNGJeblrLwIPy/aq8icxopX8mcWc=
`pragma protect end_protected
