// NIOS_test_board.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module NIOS_test_board (
		input  wire        clk_in_clk,      //    clk_in.clk
		output wire [7:0]  pio_led_export,  //   pio_led.export
		input  wire [2:0]  pio_mode_export, //  pio_mode.export
		input  wire        reset_reset_n,   //     reset.reset_n
		output wire [11:0] sdram_addr,      //     sdram.addr
		output wire [1:0]  sdram_ba,        //          .ba
		output wire        sdram_cas_n,     //          .cas_n
		output wire        sdram_cke,       //          .cke
		output wire        sdram_cs_n,      //          .cs_n
		inout  wire [15:0] sdram_dq,        //          .dq
		output wire [1:0]  sdram_dqm,       //          .dqm
		output wire        sdram_ras_n,     //          .ras_n
		output wire        sdram_we_n,      //          .we_n
		output wire        sdram_clk_clk,   // sdram_clk.clk
		input  wire        spi_g_sen_MISO,  // spi_g_sen.MISO
		output wire        spi_g_sen_MOSI,  //          .MOSI
		output wire        spi_g_sen_SCLK,  //          .SCLK
		output wire        spi_g_sen_SS_n,  //          .SS_n
		input  wire        uart_rxd,        //      uart.rxd
		output wire        uart_txd         //          .txd
	);

	wire         pll_c0_clk;                                                 // pll:c0 -> [irq_mapper:clk, mm_interconnect_0:pll_c0_clk, nios2:clk, onchip_ram:clk, pio_led:clk, pio_mode:clk, rst_controller:clk, sdram_controller:clk, spi_g_sensor:clk, sysid:clock, uart:clk]
	wire  [31:0] nios2_data_master_readdata;                                 // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                              // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                              // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [24:0] nios2_data_master_address;                                  // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                               // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                     // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                    // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                          // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                       // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [24:0] nios2_instruction_master_address;                           // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                              // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;             // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;              // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;           // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;        // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;            // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;               // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;         // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;              // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;          // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                   // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                    // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                       // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                      // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                  // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                 // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                   // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_ram_s1_address;                    // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                 // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                      // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                  // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                      // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;           // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;             // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;          // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_controller_s1_address;              // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                 // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;           // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;        // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;            // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_pio_led_s1_chipselect;                    // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                      // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                       // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                         // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                     // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                       // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                         // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                          // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                             // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                    // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                            // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                        // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire  [31:0] mm_interconnect_0_pio_mode_s1_readdata;                     // pio_mode:readdata -> mm_interconnect_0:pio_mode_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_mode_s1_address;                      // mm_interconnect_0:pio_mode_s1_address -> pio_mode:address
	wire         mm_interconnect_0_spi_g_sensor_spi_control_port_chipselect; // mm_interconnect_0:spi_g_sensor_spi_control_port_chipselect -> spi_g_sensor:spi_select
	wire  [15:0] mm_interconnect_0_spi_g_sensor_spi_control_port_readdata;   // spi_g_sensor:data_to_cpu -> mm_interconnect_0:spi_g_sensor_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_g_sensor_spi_control_port_address;    // mm_interconnect_0:spi_g_sensor_spi_control_port_address -> spi_g_sensor:mem_addr
	wire         mm_interconnect_0_spi_g_sensor_spi_control_port_read;       // mm_interconnect_0:spi_g_sensor_spi_control_port_read -> spi_g_sensor:read_n
	wire         mm_interconnect_0_spi_g_sensor_spi_control_port_write;      // mm_interconnect_0:spi_g_sensor_spi_control_port_write -> spi_g_sensor:write_n
	wire  [15:0] mm_interconnect_0_spi_g_sensor_spi_control_port_writedata;  // mm_interconnect_0:spi_g_sensor_spi_control_port_writedata -> spi_g_sensor:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                   // uart:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // spi_g_sensor:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                              // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, onchip_ram:reset, pio_led:reset_n, pio_mode:reset_n, rst_translator:in_reset, sdram_controller:reset_n, spi_g_sensor:reset_n, sysid:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                            // nios2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	NIOS_test_board_nios2 nios2 (
		.clk                                 (pll_c0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	NIOS_test_board_onchip_ram onchip_ram (
		.clk        (pll_c0_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	NIOS_test_board_pio_led pio_led (
		.clk        (pll_c0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	NIOS_test_board_pio_mode pio_mode (
		.clk      (pll_c0_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_pio_mode_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_mode_s1_readdata), //                    .readdata
		.in_port  (pio_mode_export)                         // external_connection.export
	);

	NIOS_test_board_pll pll (
		.clk                (clk_in_clk),                                //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                             //                    c1.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0)                                       //           (terminated)
	);

	NIOS_test_board_sdram_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	NIOS_test_board_spi_g_sensor spi_g_sensor (
		.clk           (pll_c0_clk),                                                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                            //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_g_sensor_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_g_sensor_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_g_sensor_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_g_sensor_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_g_sensor_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_g_sensor_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                                   //              irq.irq
		.MISO          (spi_g_sen_MISO),                                             //         external.export
		.MOSI          (spi_g_sen_MOSI),                                             //                 .export
		.SCLK          (spi_g_sen_SCLK),                                             //                 .export
		.SS_n          (spi_g_sen_SS_n)                                              //                 .export
	);

	NIOS_test_board_sysid sysid (
		.clock    (pll_c0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	NIOS_test_board_uart uart (
		.clk           (pll_c0_clk),                              //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver0_irq)                 //                 irq.irq
	);

	NIOS_test_board_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                           (clk_in_clk),                                                 //                                         clk_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                 //                                          pll_c0.clk
		.nios2_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                             //               nios2_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                             (nios2_data_master_address),                                  //                               nios2_data_master.address
		.nios2_data_master_waitrequest                         (nios2_data_master_waitrequest),                              //                                                .waitrequest
		.nios2_data_master_byteenable                          (nios2_data_master_byteenable),                               //                                                .byteenable
		.nios2_data_master_read                                (nios2_data_master_read),                                     //                                                .read
		.nios2_data_master_readdata                            (nios2_data_master_readdata),                                 //                                                .readdata
		.nios2_data_master_write                               (nios2_data_master_write),                                    //                                                .write
		.nios2_data_master_writedata                           (nios2_data_master_writedata),                                //                                                .writedata
		.nios2_data_master_debugaccess                         (nios2_data_master_debugaccess),                              //                                                .debugaccess
		.nios2_instruction_master_address                      (nios2_instruction_master_address),                           //                        nios2_instruction_master.address
		.nios2_instruction_master_waitrequest                  (nios2_instruction_master_waitrequest),                       //                                                .waitrequest
		.nios2_instruction_master_read                         (nios2_instruction_master_read),                              //                                                .read
		.nios2_instruction_master_readdata                     (nios2_instruction_master_readdata),                          //                                                .readdata
		.nios2_debug_mem_slave_address                         (mm_interconnect_0_nios2_debug_mem_slave_address),            //                           nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                           (mm_interconnect_0_nios2_debug_mem_slave_write),              //                                                .write
		.nios2_debug_mem_slave_read                            (mm_interconnect_0_nios2_debug_mem_slave_read),               //                                                .read
		.nios2_debug_mem_slave_readdata                        (mm_interconnect_0_nios2_debug_mem_slave_readdata),           //                                                .readdata
		.nios2_debug_mem_slave_writedata                       (mm_interconnect_0_nios2_debug_mem_slave_writedata),          //                                                .writedata
		.nios2_debug_mem_slave_byteenable                      (mm_interconnect_0_nios2_debug_mem_slave_byteenable),         //                                                .byteenable
		.nios2_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),        //                                                .waitrequest
		.nios2_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),        //                                                .debugaccess
		.onchip_ram_s1_address                                 (mm_interconnect_0_onchip_ram_s1_address),                    //                                   onchip_ram_s1.address
		.onchip_ram_s1_write                                   (mm_interconnect_0_onchip_ram_s1_write),                      //                                                .write
		.onchip_ram_s1_readdata                                (mm_interconnect_0_onchip_ram_s1_readdata),                   //                                                .readdata
		.onchip_ram_s1_writedata                               (mm_interconnect_0_onchip_ram_s1_writedata),                  //                                                .writedata
		.onchip_ram_s1_byteenable                              (mm_interconnect_0_onchip_ram_s1_byteenable),                 //                                                .byteenable
		.onchip_ram_s1_chipselect                              (mm_interconnect_0_onchip_ram_s1_chipselect),                 //                                                .chipselect
		.onchip_ram_s1_clken                                   (mm_interconnect_0_onchip_ram_s1_clken),                      //                                                .clken
		.pio_led_s1_address                                    (mm_interconnect_0_pio_led_s1_address),                       //                                      pio_led_s1.address
		.pio_led_s1_write                                      (mm_interconnect_0_pio_led_s1_write),                         //                                                .write
		.pio_led_s1_readdata                                   (mm_interconnect_0_pio_led_s1_readdata),                      //                                                .readdata
		.pio_led_s1_writedata                                  (mm_interconnect_0_pio_led_s1_writedata),                     //                                                .writedata
		.pio_led_s1_chipselect                                 (mm_interconnect_0_pio_led_s1_chipselect),                    //                                                .chipselect
		.pio_mode_s1_address                                   (mm_interconnect_0_pio_mode_s1_address),                      //                                     pio_mode_s1.address
		.pio_mode_s1_readdata                                  (mm_interconnect_0_pio_mode_s1_readdata),                     //                                                .readdata
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                    //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                      //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                       //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                   //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                  //                                                .writedata
		.sdram_controller_s1_address                           (mm_interconnect_0_sdram_controller_s1_address),              //                             sdram_controller_s1.address
		.sdram_controller_s1_write                             (mm_interconnect_0_sdram_controller_s1_write),                //                                                .write
		.sdram_controller_s1_read                              (mm_interconnect_0_sdram_controller_s1_read),                 //                                                .read
		.sdram_controller_s1_readdata                          (mm_interconnect_0_sdram_controller_s1_readdata),             //                                                .readdata
		.sdram_controller_s1_writedata                         (mm_interconnect_0_sdram_controller_s1_writedata),            //                                                .writedata
		.sdram_controller_s1_byteenable                        (mm_interconnect_0_sdram_controller_s1_byteenable),           //                                                .byteenable
		.sdram_controller_s1_readdatavalid                     (mm_interconnect_0_sdram_controller_s1_readdatavalid),        //                                                .readdatavalid
		.sdram_controller_s1_waitrequest                       (mm_interconnect_0_sdram_controller_s1_waitrequest),          //                                                .waitrequest
		.sdram_controller_s1_chipselect                        (mm_interconnect_0_sdram_controller_s1_chipselect),           //                                                .chipselect
		.spi_g_sensor_spi_control_port_address                 (mm_interconnect_0_spi_g_sensor_spi_control_port_address),    //                   spi_g_sensor_spi_control_port.address
		.spi_g_sensor_spi_control_port_write                   (mm_interconnect_0_spi_g_sensor_spi_control_port_write),      //                                                .write
		.spi_g_sensor_spi_control_port_read                    (mm_interconnect_0_spi_g_sensor_spi_control_port_read),       //                                                .read
		.spi_g_sensor_spi_control_port_readdata                (mm_interconnect_0_spi_g_sensor_spi_control_port_readdata),   //                                                .readdata
		.spi_g_sensor_spi_control_port_writedata               (mm_interconnect_0_spi_g_sensor_spi_control_port_writedata),  //                                                .writedata
		.spi_g_sensor_spi_control_port_chipselect              (mm_interconnect_0_spi_g_sensor_spi_control_port_chipselect), //                                                .chipselect
		.sysid_control_slave_address                           (mm_interconnect_0_sysid_control_slave_address),              //                             sysid_control_slave.address
		.sysid_control_slave_readdata                          (mm_interconnect_0_sysid_control_slave_readdata),             //                                                .readdata
		.uart_s1_address                                       (mm_interconnect_0_uart_s1_address),                          //                                         uart_s1.address
		.uart_s1_write                                         (mm_interconnect_0_uart_s1_write),                            //                                                .write
		.uart_s1_read                                          (mm_interconnect_0_uart_s1_read),                             //                                                .read
		.uart_s1_readdata                                      (mm_interconnect_0_uart_s1_readdata),                         //                                                .readdata
		.uart_s1_writedata                                     (mm_interconnect_0_uart_s1_writedata),                        //                                                .writedata
		.uart_s1_begintransfer                                 (mm_interconnect_0_uart_s1_begintransfer),                    //                                                .begintransfer
		.uart_s1_chipselect                                    (mm_interconnect_0_uart_s1_chipselect)                        //                                                .chipselect
	);

	NIOS_test_board_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_in_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
